// �Զ����ɵ�ROMģ��
// ͼƬ�ߴ�: 240 x 180
// ��ɫ��ʽ: �ڰ�(1λ)
// ���ݴ�С: 5400 �ֽ�
// ���ɹ���: image_processor.py

module Begging_240x180_rom (
    input wire clk,
    input wire [12:0] addr,
    output reg [7:0] data
);

    // ROM���ݴ洢 (5400 ����ַ)
    always @(posedge clk) begin
        case (addr)
            13'd0: data <= 8'h00;
            13'd1: data <= 8'h00;
            13'd2: data <= 8'h00;
            13'd3: data <= 8'h00;
            13'd4: data <= 8'h00;
            13'd5: data <= 8'h03;
            13'd6: data <= 8'hFF;
            13'd7: data <= 8'hFF;
            13'd8: data <= 8'hFF;
            13'd9: data <= 8'hFF;
            13'd10: data <= 8'hFF;
            13'd11: data <= 8'hFF;
            13'd12: data <= 8'hFF;
            13'd13: data <= 8'hFF;
            13'd14: data <= 8'hFF;
            13'd15: data <= 8'hFF;
            13'd16: data <= 8'hFF;
            13'd17: data <= 8'hFF;
            13'd18: data <= 8'hFF;
            13'd19: data <= 8'hFF;
            13'd20: data <= 8'hFF;
            13'd21: data <= 8'hFF;
            13'd22: data <= 8'hFF;
            13'd23: data <= 8'hFF;
            13'd24: data <= 8'h80;
            13'd25: data <= 8'h00;
            13'd26: data <= 8'h00;
            13'd27: data <= 8'h00;
            13'd28: data <= 8'h00;
            13'd29: data <= 8'h00;
            13'd30: data <= 8'h00;
            13'd31: data <= 8'h00;
            13'd32: data <= 8'h00;
            13'd33: data <= 8'h00;
            13'd34: data <= 8'h00;
            13'd35: data <= 8'h03;
            13'd36: data <= 8'hFF;
            13'd37: data <= 8'hFF;
            13'd38: data <= 8'hFF;
            13'd39: data <= 8'hFF;
            13'd40: data <= 8'hFF;
            13'd41: data <= 8'hFF;
            13'd42: data <= 8'hFF;
            13'd43: data <= 8'hFF;
            13'd44: data <= 8'hFF;
            13'd45: data <= 8'hFF;
            13'd46: data <= 8'hFF;
            13'd47: data <= 8'hFF;
            13'd48: data <= 8'hFF;
            13'd49: data <= 8'hFF;
            13'd50: data <= 8'hFF;
            13'd51: data <= 8'hFF;
            13'd52: data <= 8'hFF;
            13'd53: data <= 8'hFF;
            13'd54: data <= 8'h80;
            13'd55: data <= 8'h00;
            13'd56: data <= 8'h00;
            13'd57: data <= 8'h00;
            13'd58: data <= 8'h00;
            13'd59: data <= 8'h00;
            13'd60: data <= 8'h00;
            13'd61: data <= 8'h00;
            13'd62: data <= 8'h00;
            13'd63: data <= 8'h00;
            13'd64: data <= 8'h00;
            13'd65: data <= 8'h03;
            13'd66: data <= 8'hFF;
            13'd67: data <= 8'hFF;
            13'd68: data <= 8'hFF;
            13'd69: data <= 8'hFF;
            13'd70: data <= 8'hFF;
            13'd71: data <= 8'hFF;
            13'd72: data <= 8'hFF;
            13'd73: data <= 8'hFF;
            13'd74: data <= 8'hFF;
            13'd75: data <= 8'hFF;
            13'd76: data <= 8'hFF;
            13'd77: data <= 8'hFF;
            13'd78: data <= 8'hFF;
            13'd79: data <= 8'hFF;
            13'd80: data <= 8'hFF;
            13'd81: data <= 8'hFF;
            13'd82: data <= 8'hFF;
            13'd83: data <= 8'hFF;
            13'd84: data <= 8'h80;
            13'd85: data <= 8'h00;
            13'd86: data <= 8'h00;
            13'd87: data <= 8'h00;
            13'd88: data <= 8'h00;
            13'd89: data <= 8'h00;
            13'd90: data <= 8'h00;
            13'd91: data <= 8'h00;
            13'd92: data <= 8'h00;
            13'd93: data <= 8'h00;
            13'd94: data <= 8'h00;
            13'd95: data <= 8'h03;
            13'd96: data <= 8'hFF;
            13'd97: data <= 8'hFF;
            13'd98: data <= 8'hFF;
            13'd99: data <= 8'hFF;
            13'd100: data <= 8'hFF;
            13'd101: data <= 8'hFF;
            13'd102: data <= 8'hFF;
            13'd103: data <= 8'hFF;
            13'd104: data <= 8'hFF;
            13'd105: data <= 8'hFF;
            13'd106: data <= 8'hFF;
            13'd107: data <= 8'hFF;
            13'd108: data <= 8'hFF;
            13'd109: data <= 8'hFF;
            13'd110: data <= 8'hFF;
            13'd111: data <= 8'hFF;
            13'd112: data <= 8'hFF;
            13'd113: data <= 8'hFF;
            13'd114: data <= 8'h80;
            13'd115: data <= 8'h00;
            13'd116: data <= 8'h00;
            13'd117: data <= 8'h00;
            13'd118: data <= 8'h00;
            13'd119: data <= 8'h00;
            13'd120: data <= 8'h00;
            13'd121: data <= 8'h00;
            13'd122: data <= 8'h00;
            13'd123: data <= 8'h00;
            13'd124: data <= 8'h00;
            13'd125: data <= 8'h03;
            13'd126: data <= 8'hFF;
            13'd127: data <= 8'hFF;
            13'd128: data <= 8'hFF;
            13'd129: data <= 8'hFF;
            13'd130: data <= 8'hFF;
            13'd131: data <= 8'hFF;
            13'd132: data <= 8'hFF;
            13'd133: data <= 8'hFF;
            13'd134: data <= 8'hFF;
            13'd135: data <= 8'hFF;
            13'd136: data <= 8'hFF;
            13'd137: data <= 8'hFF;
            13'd138: data <= 8'hFF;
            13'd139: data <= 8'hFF;
            13'd140: data <= 8'hFF;
            13'd141: data <= 8'hFF;
            13'd142: data <= 8'hFF;
            13'd143: data <= 8'hFF;
            13'd144: data <= 8'h80;
            13'd145: data <= 8'h00;
            13'd146: data <= 8'h00;
            13'd147: data <= 8'h00;
            13'd148: data <= 8'h00;
            13'd149: data <= 8'h00;
            13'd150: data <= 8'h00;
            13'd151: data <= 8'h00;
            13'd152: data <= 8'h00;
            13'd153: data <= 8'h00;
            13'd154: data <= 8'h00;
            13'd155: data <= 8'h03;
            13'd156: data <= 8'hFF;
            13'd157: data <= 8'hFF;
            13'd158: data <= 8'hFF;
            13'd159: data <= 8'hFF;
            13'd160: data <= 8'hFF;
            13'd161: data <= 8'hFF;
            13'd162: data <= 8'hFF;
            13'd163: data <= 8'hFF;
            13'd164: data <= 8'hFF;
            13'd165: data <= 8'hFF;
            13'd166: data <= 8'hFF;
            13'd167: data <= 8'hFF;
            13'd168: data <= 8'hFF;
            13'd169: data <= 8'hFF;
            13'd170: data <= 8'hFF;
            13'd171: data <= 8'hFF;
            13'd172: data <= 8'hFF;
            13'd173: data <= 8'hFF;
            13'd174: data <= 8'h80;
            13'd175: data <= 8'h00;
            13'd176: data <= 8'h00;
            13'd177: data <= 8'h00;
            13'd178: data <= 8'h00;
            13'd179: data <= 8'h00;
            13'd180: data <= 8'h00;
            13'd181: data <= 8'h00;
            13'd182: data <= 8'h00;
            13'd183: data <= 8'h00;
            13'd184: data <= 8'h00;
            13'd185: data <= 8'h03;
            13'd186: data <= 8'hFF;
            13'd187: data <= 8'hFF;
            13'd188: data <= 8'hFF;
            13'd189: data <= 8'hFF;
            13'd190: data <= 8'hFF;
            13'd191: data <= 8'hFF;
            13'd192: data <= 8'hFF;
            13'd193: data <= 8'hFF;
            13'd194: data <= 8'hFF;
            13'd195: data <= 8'hFF;
            13'd196: data <= 8'hFF;
            13'd197: data <= 8'hFF;
            13'd198: data <= 8'hFF;
            13'd199: data <= 8'hFF;
            13'd200: data <= 8'hFF;
            13'd201: data <= 8'hFF;
            13'd202: data <= 8'hFF;
            13'd203: data <= 8'hFF;
            13'd204: data <= 8'h80;
            13'd205: data <= 8'h00;
            13'd206: data <= 8'h00;
            13'd207: data <= 8'h00;
            13'd208: data <= 8'h00;
            13'd209: data <= 8'h00;
            13'd210: data <= 8'h00;
            13'd211: data <= 8'h00;
            13'd212: data <= 8'h00;
            13'd213: data <= 8'h00;
            13'd214: data <= 8'h00;
            13'd215: data <= 8'h03;
            13'd216: data <= 8'hFF;
            13'd217: data <= 8'hFF;
            13'd218: data <= 8'hFF;
            13'd219: data <= 8'hFF;
            13'd220: data <= 8'hFF;
            13'd221: data <= 8'hFF;
            13'd222: data <= 8'hFF;
            13'd223: data <= 8'hFF;
            13'd224: data <= 8'hFF;
            13'd225: data <= 8'hFF;
            13'd226: data <= 8'hFF;
            13'd227: data <= 8'hFF;
            13'd228: data <= 8'hFF;
            13'd229: data <= 8'hFF;
            13'd230: data <= 8'hFF;
            13'd231: data <= 8'hFF;
            13'd232: data <= 8'hFF;
            13'd233: data <= 8'hFF;
            13'd234: data <= 8'h80;
            13'd235: data <= 8'h00;
            13'd236: data <= 8'h00;
            13'd237: data <= 8'h00;
            13'd238: data <= 8'h00;
            13'd239: data <= 8'h00;
            13'd240: data <= 8'h00;
            13'd241: data <= 8'h00;
            13'd242: data <= 8'h00;
            13'd243: data <= 8'h00;
            13'd244: data <= 8'h00;
            13'd245: data <= 8'h03;
            13'd246: data <= 8'hFF;
            13'd247: data <= 8'hFF;
            13'd248: data <= 8'hFF;
            13'd249: data <= 8'hFF;
            13'd250: data <= 8'hFF;
            13'd251: data <= 8'hFF;
            13'd252: data <= 8'hFF;
            13'd253: data <= 8'hFF;
            13'd254: data <= 8'hFF;
            13'd255: data <= 8'hFF;
            13'd256: data <= 8'hFF;
            13'd257: data <= 8'hFF;
            13'd258: data <= 8'hFF;
            13'd259: data <= 8'hFF;
            13'd260: data <= 8'hFF;
            13'd261: data <= 8'hFF;
            13'd262: data <= 8'hFF;
            13'd263: data <= 8'hFF;
            13'd264: data <= 8'h80;
            13'd265: data <= 8'h00;
            13'd266: data <= 8'h00;
            13'd267: data <= 8'h00;
            13'd268: data <= 8'h00;
            13'd269: data <= 8'h00;
            13'd270: data <= 8'h00;
            13'd271: data <= 8'h00;
            13'd272: data <= 8'h00;
            13'd273: data <= 8'h00;
            13'd274: data <= 8'h00;
            13'd275: data <= 8'h03;
            13'd276: data <= 8'hFF;
            13'd277: data <= 8'hFF;
            13'd278: data <= 8'hFF;
            13'd279: data <= 8'hFF;
            13'd280: data <= 8'hFF;
            13'd281: data <= 8'hFF;
            13'd282: data <= 8'hFF;
            13'd283: data <= 8'hFF;
            13'd284: data <= 8'hFF;
            13'd285: data <= 8'hFF;
            13'd286: data <= 8'hFF;
            13'd287: data <= 8'hFF;
            13'd288: data <= 8'hFF;
            13'd289: data <= 8'hFF;
            13'd290: data <= 8'hFF;
            13'd291: data <= 8'hFF;
            13'd292: data <= 8'hFF;
            13'd293: data <= 8'hFF;
            13'd294: data <= 8'h80;
            13'd295: data <= 8'h00;
            13'd296: data <= 8'h00;
            13'd297: data <= 8'h00;
            13'd298: data <= 8'h00;
            13'd299: data <= 8'h00;
            13'd300: data <= 8'h00;
            13'd301: data <= 8'h00;
            13'd302: data <= 8'h00;
            13'd303: data <= 8'h00;
            13'd304: data <= 8'h00;
            13'd305: data <= 8'h03;
            13'd306: data <= 8'hFF;
            13'd307: data <= 8'hFF;
            13'd308: data <= 8'hFF;
            13'd309: data <= 8'hFF;
            13'd310: data <= 8'hFF;
            13'd311: data <= 8'hFF;
            13'd312: data <= 8'hFF;
            13'd313: data <= 8'hFF;
            13'd314: data <= 8'hFF;
            13'd315: data <= 8'hFF;
            13'd316: data <= 8'hFF;
            13'd317: data <= 8'hFF;
            13'd318: data <= 8'hFF;
            13'd319: data <= 8'hFF;
            13'd320: data <= 8'hFF;
            13'd321: data <= 8'hFF;
            13'd322: data <= 8'hFF;
            13'd323: data <= 8'hFF;
            13'd324: data <= 8'h80;
            13'd325: data <= 8'h00;
            13'd326: data <= 8'h00;
            13'd327: data <= 8'h00;
            13'd328: data <= 8'h00;
            13'd329: data <= 8'h00;
            13'd330: data <= 8'h00;
            13'd331: data <= 8'h00;
            13'd332: data <= 8'h00;
            13'd333: data <= 8'h00;
            13'd334: data <= 8'h00;
            13'd335: data <= 8'h03;
            13'd336: data <= 8'hFF;
            13'd337: data <= 8'hFF;
            13'd338: data <= 8'hFF;
            13'd339: data <= 8'hFF;
            13'd340: data <= 8'hFF;
            13'd341: data <= 8'hFF;
            13'd342: data <= 8'hFF;
            13'd343: data <= 8'hFF;
            13'd344: data <= 8'hFF;
            13'd345: data <= 8'hFF;
            13'd346: data <= 8'hFF;
            13'd347: data <= 8'hFF;
            13'd348: data <= 8'hFF;
            13'd349: data <= 8'hFF;
            13'd350: data <= 8'hFF;
            13'd351: data <= 8'hFF;
            13'd352: data <= 8'hFF;
            13'd353: data <= 8'hFF;
            13'd354: data <= 8'h80;
            13'd355: data <= 8'h00;
            13'd356: data <= 8'h00;
            13'd357: data <= 8'h00;
            13'd358: data <= 8'h00;
            13'd359: data <= 8'h00;
            13'd360: data <= 8'h00;
            13'd361: data <= 8'h00;
            13'd362: data <= 8'h00;
            13'd363: data <= 8'h00;
            13'd364: data <= 8'h00;
            13'd365: data <= 8'h03;
            13'd366: data <= 8'hFF;
            13'd367: data <= 8'hFF;
            13'd368: data <= 8'hFF;
            13'd369: data <= 8'hFF;
            13'd370: data <= 8'hFF;
            13'd371: data <= 8'hFF;
            13'd372: data <= 8'hFF;
            13'd373: data <= 8'hFF;
            13'd374: data <= 8'hFF;
            13'd375: data <= 8'hFF;
            13'd376: data <= 8'hFF;
            13'd377: data <= 8'hFF;
            13'd378: data <= 8'hFF;
            13'd379: data <= 8'hFF;
            13'd380: data <= 8'hFF;
            13'd381: data <= 8'hFF;
            13'd382: data <= 8'hFF;
            13'd383: data <= 8'hFF;
            13'd384: data <= 8'h80;
            13'd385: data <= 8'h00;
            13'd386: data <= 8'h00;
            13'd387: data <= 8'h00;
            13'd388: data <= 8'h00;
            13'd389: data <= 8'h00;
            13'd390: data <= 8'h00;
            13'd391: data <= 8'h00;
            13'd392: data <= 8'h00;
            13'd393: data <= 8'h00;
            13'd394: data <= 8'h00;
            13'd395: data <= 8'h03;
            13'd396: data <= 8'hFF;
            13'd397: data <= 8'hFF;
            13'd398: data <= 8'hFF;
            13'd399: data <= 8'hFF;
            13'd400: data <= 8'hFF;
            13'd401: data <= 8'hFF;
            13'd402: data <= 8'hFF;
            13'd403: data <= 8'hFF;
            13'd404: data <= 8'hFF;
            13'd405: data <= 8'hFF;
            13'd406: data <= 8'hFF;
            13'd407: data <= 8'hFF;
            13'd408: data <= 8'hFF;
            13'd409: data <= 8'hFF;
            13'd410: data <= 8'hFF;
            13'd411: data <= 8'hFF;
            13'd412: data <= 8'hFF;
            13'd413: data <= 8'hFF;
            13'd414: data <= 8'h80;
            13'd415: data <= 8'h00;
            13'd416: data <= 8'h00;
            13'd417: data <= 8'h00;
            13'd418: data <= 8'h00;
            13'd419: data <= 8'h00;
            13'd420: data <= 8'h00;
            13'd421: data <= 8'h00;
            13'd422: data <= 8'h00;
            13'd423: data <= 8'h00;
            13'd424: data <= 8'h00;
            13'd425: data <= 8'h03;
            13'd426: data <= 8'hFF;
            13'd427: data <= 8'hFF;
            13'd428: data <= 8'hFF;
            13'd429: data <= 8'hFF;
            13'd430: data <= 8'hFF;
            13'd431: data <= 8'hFF;
            13'd432: data <= 8'hFF;
            13'd433: data <= 8'hFF;
            13'd434: data <= 8'hFF;
            13'd435: data <= 8'hFF;
            13'd436: data <= 8'hFF;
            13'd437: data <= 8'hFF;
            13'd438: data <= 8'hFF;
            13'd439: data <= 8'hFF;
            13'd440: data <= 8'hFF;
            13'd441: data <= 8'hFF;
            13'd442: data <= 8'hFF;
            13'd443: data <= 8'hFF;
            13'd444: data <= 8'h80;
            13'd445: data <= 8'h00;
            13'd446: data <= 8'h00;
            13'd447: data <= 8'h00;
            13'd448: data <= 8'h00;
            13'd449: data <= 8'h00;
            13'd450: data <= 8'h00;
            13'd451: data <= 8'h00;
            13'd452: data <= 8'h00;
            13'd453: data <= 8'h00;
            13'd454: data <= 8'h00;
            13'd455: data <= 8'h03;
            13'd456: data <= 8'hFF;
            13'd457: data <= 8'hFF;
            13'd458: data <= 8'hFF;
            13'd459: data <= 8'hFF;
            13'd460: data <= 8'hFF;
            13'd461: data <= 8'hFF;
            13'd462: data <= 8'hFF;
            13'd463: data <= 8'hFF;
            13'd464: data <= 8'hFF;
            13'd465: data <= 8'hFF;
            13'd466: data <= 8'hFF;
            13'd467: data <= 8'hFF;
            13'd468: data <= 8'hFF;
            13'd469: data <= 8'hFF;
            13'd470: data <= 8'hFF;
            13'd471: data <= 8'hFF;
            13'd472: data <= 8'hFF;
            13'd473: data <= 8'hFF;
            13'd474: data <= 8'h80;
            13'd475: data <= 8'h00;
            13'd476: data <= 8'h00;
            13'd477: data <= 8'h00;
            13'd478: data <= 8'h00;
            13'd479: data <= 8'h00;
            13'd480: data <= 8'h00;
            13'd481: data <= 8'h00;
            13'd482: data <= 8'h00;
            13'd483: data <= 8'h00;
            13'd484: data <= 8'h00;
            13'd485: data <= 8'h03;
            13'd486: data <= 8'hFF;
            13'd487: data <= 8'hFF;
            13'd488: data <= 8'hFF;
            13'd489: data <= 8'hFF;
            13'd490: data <= 8'hFF;
            13'd491: data <= 8'hFF;
            13'd492: data <= 8'hFF;
            13'd493: data <= 8'hFF;
            13'd494: data <= 8'hFF;
            13'd495: data <= 8'hFF;
            13'd496: data <= 8'hFF;
            13'd497: data <= 8'hFF;
            13'd498: data <= 8'hFF;
            13'd499: data <= 8'hFF;
            13'd500: data <= 8'hFF;
            13'd501: data <= 8'hFF;
            13'd502: data <= 8'hFF;
            13'd503: data <= 8'hFF;
            13'd504: data <= 8'h80;
            13'd505: data <= 8'h00;
            13'd506: data <= 8'h00;
            13'd507: data <= 8'h00;
            13'd508: data <= 8'h00;
            13'd509: data <= 8'h00;
            13'd510: data <= 8'h00;
            13'd511: data <= 8'h00;
            13'd512: data <= 8'h00;
            13'd513: data <= 8'h00;
            13'd514: data <= 8'h00;
            13'd515: data <= 8'h03;
            13'd516: data <= 8'hFF;
            13'd517: data <= 8'hFF;
            13'd518: data <= 8'hFF;
            13'd519: data <= 8'hFF;
            13'd520: data <= 8'hFF;
            13'd521: data <= 8'hFF;
            13'd522: data <= 8'hFF;
            13'd523: data <= 8'hFF;
            13'd524: data <= 8'hFF;
            13'd525: data <= 8'hFF;
            13'd526: data <= 8'hFF;
            13'd527: data <= 8'hFF;
            13'd528: data <= 8'hFF;
            13'd529: data <= 8'hFF;
            13'd530: data <= 8'hFF;
            13'd531: data <= 8'hFF;
            13'd532: data <= 8'hFF;
            13'd533: data <= 8'hFF;
            13'd534: data <= 8'h80;
            13'd535: data <= 8'h00;
            13'd536: data <= 8'h00;
            13'd537: data <= 8'h00;
            13'd538: data <= 8'h00;
            13'd539: data <= 8'h00;
            13'd540: data <= 8'h00;
            13'd541: data <= 8'h00;
            13'd542: data <= 8'h00;
            13'd543: data <= 8'h00;
            13'd544: data <= 8'h00;
            13'd545: data <= 8'h03;
            13'd546: data <= 8'hFF;
            13'd547: data <= 8'hFF;
            13'd548: data <= 8'hFF;
            13'd549: data <= 8'hFF;
            13'd550: data <= 8'hFF;
            13'd551: data <= 8'hFF;
            13'd552: data <= 8'hFF;
            13'd553: data <= 8'hFF;
            13'd554: data <= 8'hFF;
            13'd555: data <= 8'hFF;
            13'd556: data <= 8'hFF;
            13'd557: data <= 8'hFF;
            13'd558: data <= 8'hFF;
            13'd559: data <= 8'hFF;
            13'd560: data <= 8'hFF;
            13'd561: data <= 8'hFF;
            13'd562: data <= 8'hFF;
            13'd563: data <= 8'hFF;
            13'd564: data <= 8'h80;
            13'd565: data <= 8'h00;
            13'd566: data <= 8'h00;
            13'd567: data <= 8'h00;
            13'd568: data <= 8'h00;
            13'd569: data <= 8'h00;
            13'd570: data <= 8'h00;
            13'd571: data <= 8'h00;
            13'd572: data <= 8'h00;
            13'd573: data <= 8'h00;
            13'd574: data <= 8'h00;
            13'd575: data <= 8'h03;
            13'd576: data <= 8'hFF;
            13'd577: data <= 8'hFF;
            13'd578: data <= 8'hFF;
            13'd579: data <= 8'hFF;
            13'd580: data <= 8'hFF;
            13'd581: data <= 8'hFF;
            13'd582: data <= 8'hFF;
            13'd583: data <= 8'hFF;
            13'd584: data <= 8'hFF;
            13'd585: data <= 8'hFF;
            13'd586: data <= 8'hFF;
            13'd587: data <= 8'hFF;
            13'd588: data <= 8'hFF;
            13'd589: data <= 8'hFF;
            13'd590: data <= 8'hFF;
            13'd591: data <= 8'hFF;
            13'd592: data <= 8'hFF;
            13'd593: data <= 8'hFF;
            13'd594: data <= 8'h80;
            13'd595: data <= 8'h00;
            13'd596: data <= 8'h00;
            13'd597: data <= 8'h00;
            13'd598: data <= 8'h00;
            13'd599: data <= 8'h00;
            13'd600: data <= 8'h00;
            13'd601: data <= 8'h00;
            13'd602: data <= 8'h00;
            13'd603: data <= 8'h00;
            13'd604: data <= 8'h00;
            13'd605: data <= 8'h03;
            13'd606: data <= 8'hFF;
            13'd607: data <= 8'hFF;
            13'd608: data <= 8'hFF;
            13'd609: data <= 8'hFF;
            13'd610: data <= 8'hFF;
            13'd611: data <= 8'hFF;
            13'd612: data <= 8'hFF;
            13'd613: data <= 8'hFF;
            13'd614: data <= 8'hFF;
            13'd615: data <= 8'hFF;
            13'd616: data <= 8'hFF;
            13'd617: data <= 8'hFF;
            13'd618: data <= 8'hFF;
            13'd619: data <= 8'hFF;
            13'd620: data <= 8'hFF;
            13'd621: data <= 8'hFF;
            13'd622: data <= 8'hFF;
            13'd623: data <= 8'hFF;
            13'd624: data <= 8'h80;
            13'd625: data <= 8'h00;
            13'd626: data <= 8'h00;
            13'd627: data <= 8'h00;
            13'd628: data <= 8'h00;
            13'd629: data <= 8'h00;
            13'd630: data <= 8'h00;
            13'd631: data <= 8'h00;
            13'd632: data <= 8'h00;
            13'd633: data <= 8'h00;
            13'd634: data <= 8'h00;
            13'd635: data <= 8'h03;
            13'd636: data <= 8'hFF;
            13'd637: data <= 8'hFF;
            13'd638: data <= 8'hFF;
            13'd639: data <= 8'hFF;
            13'd640: data <= 8'hFF;
            13'd641: data <= 8'hFF;
            13'd642: data <= 8'hFF;
            13'd643: data <= 8'hFF;
            13'd644: data <= 8'hFF;
            13'd645: data <= 8'hFF;
            13'd646: data <= 8'hFF;
            13'd647: data <= 8'hFF;
            13'd648: data <= 8'hFF;
            13'd649: data <= 8'hFF;
            13'd650: data <= 8'hFF;
            13'd651: data <= 8'hFF;
            13'd652: data <= 8'hFF;
            13'd653: data <= 8'hFF;
            13'd654: data <= 8'h80;
            13'd655: data <= 8'h00;
            13'd656: data <= 8'h00;
            13'd657: data <= 8'h00;
            13'd658: data <= 8'h00;
            13'd659: data <= 8'h00;
            13'd660: data <= 8'h00;
            13'd661: data <= 8'h00;
            13'd662: data <= 8'h00;
            13'd663: data <= 8'h00;
            13'd664: data <= 8'h00;
            13'd665: data <= 8'h03;
            13'd666: data <= 8'hFF;
            13'd667: data <= 8'hFF;
            13'd668: data <= 8'hFF;
            13'd669: data <= 8'hFF;
            13'd670: data <= 8'hFF;
            13'd671: data <= 8'hFF;
            13'd672: data <= 8'hFF;
            13'd673: data <= 8'hFF;
            13'd674: data <= 8'hFF;
            13'd675: data <= 8'hFF;
            13'd676: data <= 8'hFF;
            13'd677: data <= 8'hFF;
            13'd678: data <= 8'hFF;
            13'd679: data <= 8'hFF;
            13'd680: data <= 8'hFF;
            13'd681: data <= 8'hFF;
            13'd682: data <= 8'hFF;
            13'd683: data <= 8'hFF;
            13'd684: data <= 8'h80;
            13'd685: data <= 8'h00;
            13'd686: data <= 8'h00;
            13'd687: data <= 8'h00;
            13'd688: data <= 8'h00;
            13'd689: data <= 8'h00;
            13'd690: data <= 8'h00;
            13'd691: data <= 8'h00;
            13'd692: data <= 8'h00;
            13'd693: data <= 8'h00;
            13'd694: data <= 8'h00;
            13'd695: data <= 8'h03;
            13'd696: data <= 8'hFF;
            13'd697: data <= 8'hFF;
            13'd698: data <= 8'hFF;
            13'd699: data <= 8'hFF;
            13'd700: data <= 8'hFF;
            13'd701: data <= 8'hFF;
            13'd702: data <= 8'hFF;
            13'd703: data <= 8'hFF;
            13'd704: data <= 8'hFF;
            13'd705: data <= 8'hFF;
            13'd706: data <= 8'hFF;
            13'd707: data <= 8'hFF;
            13'd708: data <= 8'hFF;
            13'd709: data <= 8'hFF;
            13'd710: data <= 8'hFF;
            13'd711: data <= 8'hFF;
            13'd712: data <= 8'hFF;
            13'd713: data <= 8'hFF;
            13'd714: data <= 8'h80;
            13'd715: data <= 8'h00;
            13'd716: data <= 8'h00;
            13'd717: data <= 8'h00;
            13'd718: data <= 8'h00;
            13'd719: data <= 8'h00;
            13'd720: data <= 8'h00;
            13'd721: data <= 8'h00;
            13'd722: data <= 8'h00;
            13'd723: data <= 8'h00;
            13'd724: data <= 8'h00;
            13'd725: data <= 8'h03;
            13'd726: data <= 8'hFF;
            13'd727: data <= 8'hFF;
            13'd728: data <= 8'hFF;
            13'd729: data <= 8'hFF;
            13'd730: data <= 8'hFF;
            13'd731: data <= 8'hFF;
            13'd732: data <= 8'hFF;
            13'd733: data <= 8'hFF;
            13'd734: data <= 8'hFF;
            13'd735: data <= 8'hFF;
            13'd736: data <= 8'hFF;
            13'd737: data <= 8'hFF;
            13'd738: data <= 8'hFF;
            13'd739: data <= 8'hFF;
            13'd740: data <= 8'hFF;
            13'd741: data <= 8'hFF;
            13'd742: data <= 8'hFF;
            13'd743: data <= 8'hFF;
            13'd744: data <= 8'h80;
            13'd745: data <= 8'h00;
            13'd746: data <= 8'h00;
            13'd747: data <= 8'h00;
            13'd748: data <= 8'h00;
            13'd749: data <= 8'h00;
            13'd750: data <= 8'h00;
            13'd751: data <= 8'h00;
            13'd752: data <= 8'h00;
            13'd753: data <= 8'h00;
            13'd754: data <= 8'h00;
            13'd755: data <= 8'h03;
            13'd756: data <= 8'hFF;
            13'd757: data <= 8'hFF;
            13'd758: data <= 8'hFF;
            13'd759: data <= 8'hFF;
            13'd760: data <= 8'hFF;
            13'd761: data <= 8'hFF;
            13'd762: data <= 8'hFF;
            13'd763: data <= 8'hFF;
            13'd764: data <= 8'hFF;
            13'd765: data <= 8'hFF;
            13'd766: data <= 8'hFF;
            13'd767: data <= 8'hFF;
            13'd768: data <= 8'hFF;
            13'd769: data <= 8'hFF;
            13'd770: data <= 8'hFF;
            13'd771: data <= 8'hFF;
            13'd772: data <= 8'hFF;
            13'd773: data <= 8'hFF;
            13'd774: data <= 8'h80;
            13'd775: data <= 8'h00;
            13'd776: data <= 8'h00;
            13'd777: data <= 8'h00;
            13'd778: data <= 8'h00;
            13'd779: data <= 8'h00;
            13'd780: data <= 8'h00;
            13'd781: data <= 8'h00;
            13'd782: data <= 8'h00;
            13'd783: data <= 8'h00;
            13'd784: data <= 8'h00;
            13'd785: data <= 8'h03;
            13'd786: data <= 8'hFF;
            13'd787: data <= 8'hFF;
            13'd788: data <= 8'hFF;
            13'd789: data <= 8'hFF;
            13'd790: data <= 8'hFF;
            13'd791: data <= 8'hFF;
            13'd792: data <= 8'hFF;
            13'd793: data <= 8'hFF;
            13'd794: data <= 8'hFF;
            13'd795: data <= 8'hFF;
            13'd796: data <= 8'hFF;
            13'd797: data <= 8'hFF;
            13'd798: data <= 8'hFF;
            13'd799: data <= 8'hFF;
            13'd800: data <= 8'hFF;
            13'd801: data <= 8'hFF;
            13'd802: data <= 8'hFF;
            13'd803: data <= 8'hFF;
            13'd804: data <= 8'h80;
            13'd805: data <= 8'h00;
            13'd806: data <= 8'h00;
            13'd807: data <= 8'h00;
            13'd808: data <= 8'h00;
            13'd809: data <= 8'h00;
            13'd810: data <= 8'h00;
            13'd811: data <= 8'h00;
            13'd812: data <= 8'h00;
            13'd813: data <= 8'h00;
            13'd814: data <= 8'h00;
            13'd815: data <= 8'h03;
            13'd816: data <= 8'hFF;
            13'd817: data <= 8'hFF;
            13'd818: data <= 8'hFF;
            13'd819: data <= 8'hFF;
            13'd820: data <= 8'hFF;
            13'd821: data <= 8'hFF;
            13'd822: data <= 8'hFF;
            13'd823: data <= 8'hFF;
            13'd824: data <= 8'hFF;
            13'd825: data <= 8'hFF;
            13'd826: data <= 8'hFF;
            13'd827: data <= 8'hFF;
            13'd828: data <= 8'hFF;
            13'd829: data <= 8'hFF;
            13'd830: data <= 8'hFF;
            13'd831: data <= 8'hFF;
            13'd832: data <= 8'hFF;
            13'd833: data <= 8'hFF;
            13'd834: data <= 8'h80;
            13'd835: data <= 8'h00;
            13'd836: data <= 8'h00;
            13'd837: data <= 8'h00;
            13'd838: data <= 8'h00;
            13'd839: data <= 8'h00;
            13'd840: data <= 8'h00;
            13'd841: data <= 8'h00;
            13'd842: data <= 8'h00;
            13'd843: data <= 8'h00;
            13'd844: data <= 8'h00;
            13'd845: data <= 8'h03;
            13'd846: data <= 8'hFF;
            13'd847: data <= 8'hFF;
            13'd848: data <= 8'hFF;
            13'd849: data <= 8'hFF;
            13'd850: data <= 8'hFF;
            13'd851: data <= 8'hFF;
            13'd852: data <= 8'hFF;
            13'd853: data <= 8'hFF;
            13'd854: data <= 8'hFF;
            13'd855: data <= 8'hFF;
            13'd856: data <= 8'hFF;
            13'd857: data <= 8'hFF;
            13'd858: data <= 8'hFF;
            13'd859: data <= 8'hFF;
            13'd860: data <= 8'hFF;
            13'd861: data <= 8'hFF;
            13'd862: data <= 8'hFF;
            13'd863: data <= 8'hFF;
            13'd864: data <= 8'h80;
            13'd865: data <= 8'h00;
            13'd866: data <= 8'h00;
            13'd867: data <= 8'h00;
            13'd868: data <= 8'h00;
            13'd869: data <= 8'h00;
            13'd870: data <= 8'h00;
            13'd871: data <= 8'h00;
            13'd872: data <= 8'h00;
            13'd873: data <= 8'h00;
            13'd874: data <= 8'h00;
            13'd875: data <= 8'h03;
            13'd876: data <= 8'hFF;
            13'd877: data <= 8'hFF;
            13'd878: data <= 8'hFF;
            13'd879: data <= 8'hFF;
            13'd880: data <= 8'hFF;
            13'd881: data <= 8'hFF;
            13'd882: data <= 8'hFF;
            13'd883: data <= 8'hFF;
            13'd884: data <= 8'hFF;
            13'd885: data <= 8'hFF;
            13'd886: data <= 8'hFF;
            13'd887: data <= 8'hFF;
            13'd888: data <= 8'hFF;
            13'd889: data <= 8'hFF;
            13'd890: data <= 8'hFF;
            13'd891: data <= 8'hFF;
            13'd892: data <= 8'hFF;
            13'd893: data <= 8'hFF;
            13'd894: data <= 8'h80;
            13'd895: data <= 8'h00;
            13'd896: data <= 8'h00;
            13'd897: data <= 8'h00;
            13'd898: data <= 8'h00;
            13'd899: data <= 8'h00;
            13'd900: data <= 8'h00;
            13'd901: data <= 8'h00;
            13'd902: data <= 8'h00;
            13'd903: data <= 8'h00;
            13'd904: data <= 8'h00;
            13'd905: data <= 8'h03;
            13'd906: data <= 8'hFF;
            13'd907: data <= 8'hFF;
            13'd908: data <= 8'hFF;
            13'd909: data <= 8'hFF;
            13'd910: data <= 8'hFF;
            13'd911: data <= 8'hFF;
            13'd912: data <= 8'hFF;
            13'd913: data <= 8'hFF;
            13'd914: data <= 8'hFF;
            13'd915: data <= 8'hE0;
            13'd916: data <= 8'hFF;
            13'd917: data <= 8'hFF;
            13'd918: data <= 8'hFF;
            13'd919: data <= 8'hFF;
            13'd920: data <= 8'hFF;
            13'd921: data <= 8'hFF;
            13'd922: data <= 8'hFF;
            13'd923: data <= 8'hFF;
            13'd924: data <= 8'h80;
            13'd925: data <= 8'h00;
            13'd926: data <= 8'h00;
            13'd927: data <= 8'h00;
            13'd928: data <= 8'h00;
            13'd929: data <= 8'h00;
            13'd930: data <= 8'h00;
            13'd931: data <= 8'h00;
            13'd932: data <= 8'h00;
            13'd933: data <= 8'h00;
            13'd934: data <= 8'h00;
            13'd935: data <= 8'h03;
            13'd936: data <= 8'hFF;
            13'd937: data <= 8'hFF;
            13'd938: data <= 8'hFF;
            13'd939: data <= 8'hFF;
            13'd940: data <= 8'hFF;
            13'd941: data <= 8'hFF;
            13'd942: data <= 8'hFF;
            13'd943: data <= 8'hFF;
            13'd944: data <= 8'hFF;
            13'd945: data <= 8'h80;
            13'd946: data <= 8'h3F;
            13'd947: data <= 8'hFF;
            13'd948: data <= 8'hFF;
            13'd949: data <= 8'hFF;
            13'd950: data <= 8'hFF;
            13'd951: data <= 8'hFF;
            13'd952: data <= 8'hFF;
            13'd953: data <= 8'hFF;
            13'd954: data <= 8'h80;
            13'd955: data <= 8'h00;
            13'd956: data <= 8'h00;
            13'd957: data <= 8'h00;
            13'd958: data <= 8'h00;
            13'd959: data <= 8'h00;
            13'd960: data <= 8'h00;
            13'd961: data <= 8'h00;
            13'd962: data <= 8'h00;
            13'd963: data <= 8'h00;
            13'd964: data <= 8'h00;
            13'd965: data <= 8'h03;
            13'd966: data <= 8'hFF;
            13'd967: data <= 8'hFF;
            13'd968: data <= 8'hFF;
            13'd969: data <= 8'hFF;
            13'd970: data <= 8'hFF;
            13'd971: data <= 8'hFF;
            13'd972: data <= 8'hFF;
            13'd973: data <= 8'hFF;
            13'd974: data <= 8'h80;
            13'd975: data <= 8'h00;
            13'd976: data <= 8'h1F;
            13'd977: data <= 8'hFF;
            13'd978: data <= 8'hFF;
            13'd979: data <= 8'hFF;
            13'd980: data <= 8'hFF;
            13'd981: data <= 8'hFF;
            13'd982: data <= 8'hFF;
            13'd983: data <= 8'hFF;
            13'd984: data <= 8'h80;
            13'd985: data <= 8'h00;
            13'd986: data <= 8'h00;
            13'd987: data <= 8'h00;
            13'd988: data <= 8'h00;
            13'd989: data <= 8'h00;
            13'd990: data <= 8'h00;
            13'd991: data <= 8'h00;
            13'd992: data <= 8'h00;
            13'd993: data <= 8'h00;
            13'd994: data <= 8'h00;
            13'd995: data <= 8'h03;
            13'd996: data <= 8'hFF;
            13'd997: data <= 8'hFF;
            13'd998: data <= 8'hFF;
            13'd999: data <= 8'hFF;
            13'd1000: data <= 8'hFF;
            13'd1001: data <= 8'hFF;
            13'd1002: data <= 8'hFF;
            13'd1003: data <= 8'h80;
            13'd1004: data <= 8'h00;
            13'd1005: data <= 8'h00;
            13'd1006: data <= 8'h1F;
            13'd1007: data <= 8'hFF;
            13'd1008: data <= 8'hFF;
            13'd1009: data <= 8'hFF;
            13'd1010: data <= 8'hFF;
            13'd1011: data <= 8'hFF;
            13'd1012: data <= 8'hFF;
            13'd1013: data <= 8'hFF;
            13'd1014: data <= 8'h80;
            13'd1015: data <= 8'h00;
            13'd1016: data <= 8'h00;
            13'd1017: data <= 8'h00;
            13'd1018: data <= 8'h00;
            13'd1019: data <= 8'h00;
            13'd1020: data <= 8'h00;
            13'd1021: data <= 8'h00;
            13'd1022: data <= 8'h00;
            13'd1023: data <= 8'h00;
            13'd1024: data <= 8'h00;
            13'd1025: data <= 8'h03;
            13'd1026: data <= 8'hFF;
            13'd1027: data <= 8'hFF;
            13'd1028: data <= 8'hFF;
            13'd1029: data <= 8'hFF;
            13'd1030: data <= 8'hFF;
            13'd1031: data <= 8'hFF;
            13'd1032: data <= 8'hFE;
            13'd1033: data <= 8'h00;
            13'd1034: data <= 8'h00;
            13'd1035: data <= 8'h00;
            13'd1036: data <= 8'h1F;
            13'd1037: data <= 8'hFF;
            13'd1038: data <= 8'hFF;
            13'd1039: data <= 8'hFF;
            13'd1040: data <= 8'hFF;
            13'd1041: data <= 8'hFF;
            13'd1042: data <= 8'hFF;
            13'd1043: data <= 8'hFF;
            13'd1044: data <= 8'h80;
            13'd1045: data <= 8'h00;
            13'd1046: data <= 8'h00;
            13'd1047: data <= 8'h00;
            13'd1048: data <= 8'h00;
            13'd1049: data <= 8'h00;
            13'd1050: data <= 8'h00;
            13'd1051: data <= 8'h00;
            13'd1052: data <= 8'h00;
            13'd1053: data <= 8'h00;
            13'd1054: data <= 8'h00;
            13'd1055: data <= 8'h03;
            13'd1056: data <= 8'hFF;
            13'd1057: data <= 8'hFF;
            13'd1058: data <= 8'hFF;
            13'd1059: data <= 8'hFF;
            13'd1060: data <= 8'hFF;
            13'd1061: data <= 8'hFF;
            13'd1062: data <= 8'h80;
            13'd1063: data <= 8'h00;
            13'd1064: data <= 8'h00;
            13'd1065: data <= 8'h00;
            13'd1066: data <= 8'h0F;
            13'd1067: data <= 8'hFF;
            13'd1068: data <= 8'hFF;
            13'd1069: data <= 8'hFF;
            13'd1070: data <= 8'hFF;
            13'd1071: data <= 8'hFF;
            13'd1072: data <= 8'hFF;
            13'd1073: data <= 8'hFF;
            13'd1074: data <= 8'h80;
            13'd1075: data <= 8'h00;
            13'd1076: data <= 8'h00;
            13'd1077: data <= 8'h00;
            13'd1078: data <= 8'h00;
            13'd1079: data <= 8'h00;
            13'd1080: data <= 8'h00;
            13'd1081: data <= 8'h00;
            13'd1082: data <= 8'h00;
            13'd1083: data <= 8'h00;
            13'd1084: data <= 8'h00;
            13'd1085: data <= 8'h03;
            13'd1086: data <= 8'hFF;
            13'd1087: data <= 8'hFF;
            13'd1088: data <= 8'hFF;
            13'd1089: data <= 8'hFF;
            13'd1090: data <= 8'hFF;
            13'd1091: data <= 8'hFE;
            13'd1092: data <= 8'h00;
            13'd1093: data <= 8'h00;
            13'd1094: data <= 8'h00;
            13'd1095: data <= 8'h00;
            13'd1096: data <= 8'h07;
            13'd1097: data <= 8'hFF;
            13'd1098: data <= 8'hFF;
            13'd1099: data <= 8'hFF;
            13'd1100: data <= 8'hFF;
            13'd1101: data <= 8'hFF;
            13'd1102: data <= 8'hFF;
            13'd1103: data <= 8'hFF;
            13'd1104: data <= 8'h80;
            13'd1105: data <= 8'h00;
            13'd1106: data <= 8'h00;
            13'd1107: data <= 8'h00;
            13'd1108: data <= 8'h00;
            13'd1109: data <= 8'h00;
            13'd1110: data <= 8'h00;
            13'd1111: data <= 8'h00;
            13'd1112: data <= 8'h00;
            13'd1113: data <= 8'h00;
            13'd1114: data <= 8'h00;
            13'd1115: data <= 8'h03;
            13'd1116: data <= 8'hFF;
            13'd1117: data <= 8'hFF;
            13'd1118: data <= 8'hFF;
            13'd1119: data <= 8'hFF;
            13'd1120: data <= 8'hFF;
            13'd1121: data <= 8'hF0;
            13'd1122: data <= 8'h00;
            13'd1123: data <= 8'h00;
            13'd1124: data <= 8'h00;
            13'd1125: data <= 8'h10;
            13'd1126: data <= 8'h07;
            13'd1127: data <= 8'hFF;
            13'd1128: data <= 8'hFF;
            13'd1129: data <= 8'hFF;
            13'd1130: data <= 8'hFF;
            13'd1131: data <= 8'hFF;
            13'd1132: data <= 8'hFF;
            13'd1133: data <= 8'hFF;
            13'd1134: data <= 8'h80;
            13'd1135: data <= 8'h00;
            13'd1136: data <= 8'h00;
            13'd1137: data <= 8'h00;
            13'd1138: data <= 8'h00;
            13'd1139: data <= 8'h00;
            13'd1140: data <= 8'h00;
            13'd1141: data <= 8'h00;
            13'd1142: data <= 8'h00;
            13'd1143: data <= 8'h00;
            13'd1144: data <= 8'h00;
            13'd1145: data <= 8'h03;
            13'd1146: data <= 8'hFF;
            13'd1147: data <= 8'hFF;
            13'd1148: data <= 8'hFF;
            13'd1149: data <= 8'hFF;
            13'd1150: data <= 8'hFF;
            13'd1151: data <= 8'hC0;
            13'd1152: data <= 8'h00;
            13'd1153: data <= 8'h00;
            13'd1154: data <= 8'h01;
            13'd1155: data <= 8'hFC;
            13'd1156: data <= 8'h03;
            13'd1157: data <= 8'hFF;
            13'd1158: data <= 8'hFF;
            13'd1159: data <= 8'hFF;
            13'd1160: data <= 8'hFF;
            13'd1161: data <= 8'hFF;
            13'd1162: data <= 8'hFF;
            13'd1163: data <= 8'hFF;
            13'd1164: data <= 8'h80;
            13'd1165: data <= 8'h00;
            13'd1166: data <= 8'h00;
            13'd1167: data <= 8'h00;
            13'd1168: data <= 8'h00;
            13'd1169: data <= 8'h00;
            13'd1170: data <= 8'h00;
            13'd1171: data <= 8'h00;
            13'd1172: data <= 8'h00;
            13'd1173: data <= 8'h00;
            13'd1174: data <= 8'h00;
            13'd1175: data <= 8'h03;
            13'd1176: data <= 8'hFF;
            13'd1177: data <= 8'hFF;
            13'd1178: data <= 8'hFF;
            13'd1179: data <= 8'hFF;
            13'd1180: data <= 8'hFE;
            13'd1181: data <= 8'h00;
            13'd1182: data <= 8'h00;
            13'd1183: data <= 8'h00;
            13'd1184: data <= 8'hFF;
            13'd1185: data <= 8'hFE;
            13'd1186: data <= 8'h00;
            13'd1187: data <= 8'h7F;
            13'd1188: data <= 8'hFF;
            13'd1189: data <= 8'hFF;
            13'd1190: data <= 8'hFF;
            13'd1191: data <= 8'hFF;
            13'd1192: data <= 8'hFF;
            13'd1193: data <= 8'hFF;
            13'd1194: data <= 8'h80;
            13'd1195: data <= 8'h00;
            13'd1196: data <= 8'h00;
            13'd1197: data <= 8'h00;
            13'd1198: data <= 8'h00;
            13'd1199: data <= 8'h00;
            13'd1200: data <= 8'h00;
            13'd1201: data <= 8'h00;
            13'd1202: data <= 8'h00;
            13'd1203: data <= 8'h00;
            13'd1204: data <= 8'h00;
            13'd1205: data <= 8'h03;
            13'd1206: data <= 8'hFF;
            13'd1207: data <= 8'hFF;
            13'd1208: data <= 8'hFF;
            13'd1209: data <= 8'hFF;
            13'd1210: data <= 8'hF8;
            13'd1211: data <= 8'h00;
            13'd1212: data <= 8'h00;
            13'd1213: data <= 8'h3F;
            13'd1214: data <= 8'hFF;
            13'd1215: data <= 8'hFE;
            13'd1216: data <= 8'h00;
            13'd1217: data <= 8'h1F;
            13'd1218: data <= 8'hFF;
            13'd1219: data <= 8'hFF;
            13'd1220: data <= 8'hFF;
            13'd1221: data <= 8'hFF;
            13'd1222: data <= 8'hFF;
            13'd1223: data <= 8'hFF;
            13'd1224: data <= 8'h80;
            13'd1225: data <= 8'h00;
            13'd1226: data <= 8'h00;
            13'd1227: data <= 8'h00;
            13'd1228: data <= 8'h00;
            13'd1229: data <= 8'h00;
            13'd1230: data <= 8'h00;
            13'd1231: data <= 8'h00;
            13'd1232: data <= 8'h00;
            13'd1233: data <= 8'h00;
            13'd1234: data <= 8'h00;
            13'd1235: data <= 8'h03;
            13'd1236: data <= 8'hFF;
            13'd1237: data <= 8'hFF;
            13'd1238: data <= 8'hFF;
            13'd1239: data <= 8'hFF;
            13'd1240: data <= 8'hC0;
            13'd1241: data <= 8'h00;
            13'd1242: data <= 8'h07;
            13'd1243: data <= 8'hFF;
            13'd1244: data <= 8'hFF;
            13'd1245: data <= 8'hFF;
            13'd1246: data <= 8'h00;
            13'd1247: data <= 8'h03;
            13'd1248: data <= 8'hFF;
            13'd1249: data <= 8'hFF;
            13'd1250: data <= 8'hFF;
            13'd1251: data <= 8'hFF;
            13'd1252: data <= 8'hFF;
            13'd1253: data <= 8'hFF;
            13'd1254: data <= 8'h80;
            13'd1255: data <= 8'h00;
            13'd1256: data <= 8'h00;
            13'd1257: data <= 8'h00;
            13'd1258: data <= 8'h00;
            13'd1259: data <= 8'h00;
            13'd1260: data <= 8'h00;
            13'd1261: data <= 8'h00;
            13'd1262: data <= 8'h00;
            13'd1263: data <= 8'h00;
            13'd1264: data <= 8'h00;
            13'd1265: data <= 8'h03;
            13'd1266: data <= 8'hFF;
            13'd1267: data <= 8'hFF;
            13'd1268: data <= 8'hFF;
            13'd1269: data <= 8'hFF;
            13'd1270: data <= 8'h00;
            13'd1271: data <= 8'h00;
            13'd1272: data <= 8'h3F;
            13'd1273: data <= 8'hFF;
            13'd1274: data <= 8'hFF;
            13'd1275: data <= 8'hFF;
            13'd1276: data <= 8'h80;
            13'd1277: data <= 8'h00;
            13'd1278: data <= 8'h7F;
            13'd1279: data <= 8'hFF;
            13'd1280: data <= 8'hFF;
            13'd1281: data <= 8'hFF;
            13'd1282: data <= 8'hFF;
            13'd1283: data <= 8'hFF;
            13'd1284: data <= 8'h80;
            13'd1285: data <= 8'h00;
            13'd1286: data <= 8'h00;
            13'd1287: data <= 8'h00;
            13'd1288: data <= 8'h00;
            13'd1289: data <= 8'h00;
            13'd1290: data <= 8'h00;
            13'd1291: data <= 8'h00;
            13'd1292: data <= 8'h00;
            13'd1293: data <= 8'h00;
            13'd1294: data <= 8'h00;
            13'd1295: data <= 8'h03;
            13'd1296: data <= 8'hFF;
            13'd1297: data <= 8'hFF;
            13'd1298: data <= 8'hFF;
            13'd1299: data <= 8'hFE;
            13'd1300: data <= 8'h00;
            13'd1301: data <= 8'h01;
            13'd1302: data <= 8'hFF;
            13'd1303: data <= 8'hFF;
            13'd1304: data <= 8'hFF;
            13'd1305: data <= 8'hFF;
            13'd1306: data <= 8'hC0;
            13'd1307: data <= 8'h00;
            13'd1308: data <= 8'h04;
            13'd1309: data <= 8'h03;
            13'd1310: data <= 8'hFF;
            13'd1311: data <= 8'hFF;
            13'd1312: data <= 8'hFF;
            13'd1313: data <= 8'hFF;
            13'd1314: data <= 8'h80;
            13'd1315: data <= 8'h00;
            13'd1316: data <= 8'h00;
            13'd1317: data <= 8'h00;
            13'd1318: data <= 8'h00;
            13'd1319: data <= 8'h00;
            13'd1320: data <= 8'h00;
            13'd1321: data <= 8'h00;
            13'd1322: data <= 8'h00;
            13'd1323: data <= 8'h00;
            13'd1324: data <= 8'h00;
            13'd1325: data <= 8'h03;
            13'd1326: data <= 8'hFF;
            13'd1327: data <= 8'hFF;
            13'd1328: data <= 8'hFF;
            13'd1329: data <= 8'hFC;
            13'd1330: data <= 8'h00;
            13'd1331: data <= 8'h0F;
            13'd1332: data <= 8'hFF;
            13'd1333: data <= 8'hFF;
            13'd1334: data <= 8'hFF;
            13'd1335: data <= 8'hFF;
            13'd1336: data <= 8'hF0;
            13'd1337: data <= 8'h00;
            13'd1338: data <= 8'h00;
            13'd1339: data <= 8'h01;
            13'd1340: data <= 8'hFF;
            13'd1341: data <= 8'hFF;
            13'd1342: data <= 8'hFF;
            13'd1343: data <= 8'hFF;
            13'd1344: data <= 8'h80;
            13'd1345: data <= 8'h00;
            13'd1346: data <= 8'h00;
            13'd1347: data <= 8'h00;
            13'd1348: data <= 8'h00;
            13'd1349: data <= 8'h00;
            13'd1350: data <= 8'h00;
            13'd1351: data <= 8'h00;
            13'd1352: data <= 8'h00;
            13'd1353: data <= 8'h00;
            13'd1354: data <= 8'h00;
            13'd1355: data <= 8'h03;
            13'd1356: data <= 8'hFF;
            13'd1357: data <= 8'hFF;
            13'd1358: data <= 8'hFF;
            13'd1359: data <= 8'hF0;
            13'd1360: data <= 8'h00;
            13'd1361: data <= 8'h7F;
            13'd1362: data <= 8'hFF;
            13'd1363: data <= 8'hFF;
            13'd1364: data <= 8'hFF;
            13'd1365: data <= 8'hFF;
            13'd1366: data <= 8'hFC;
            13'd1367: data <= 8'h00;
            13'd1368: data <= 8'h00;
            13'd1369: data <= 8'h00;
            13'd1370: data <= 8'hFF;
            13'd1371: data <= 8'hFF;
            13'd1372: data <= 8'hFF;
            13'd1373: data <= 8'hFF;
            13'd1374: data <= 8'h80;
            13'd1375: data <= 8'h00;
            13'd1376: data <= 8'h00;
            13'd1377: data <= 8'h00;
            13'd1378: data <= 8'h00;
            13'd1379: data <= 8'h00;
            13'd1380: data <= 8'h00;
            13'd1381: data <= 8'h00;
            13'd1382: data <= 8'h00;
            13'd1383: data <= 8'h00;
            13'd1384: data <= 8'h00;
            13'd1385: data <= 8'h03;
            13'd1386: data <= 8'hFF;
            13'd1387: data <= 8'hFF;
            13'd1388: data <= 8'hFF;
            13'd1389: data <= 8'hE0;
            13'd1390: data <= 8'h03;
            13'd1391: data <= 8'hFF;
            13'd1392: data <= 8'hFF;
            13'd1393: data <= 8'hFF;
            13'd1394: data <= 8'hFF;
            13'd1395: data <= 8'hFF;
            13'd1396: data <= 8'hFF;
            13'd1397: data <= 8'h00;
            13'd1398: data <= 8'h00;
            13'd1399: data <= 8'h00;
            13'd1400: data <= 8'h7F;
            13'd1401: data <= 8'hFF;
            13'd1402: data <= 8'hFF;
            13'd1403: data <= 8'hFF;
            13'd1404: data <= 8'h80;
            13'd1405: data <= 8'h00;
            13'd1406: data <= 8'h00;
            13'd1407: data <= 8'h00;
            13'd1408: data <= 8'h00;
            13'd1409: data <= 8'h00;
            13'd1410: data <= 8'h00;
            13'd1411: data <= 8'h00;
            13'd1412: data <= 8'h00;
            13'd1413: data <= 8'h00;
            13'd1414: data <= 8'h00;
            13'd1415: data <= 8'h03;
            13'd1416: data <= 8'hFF;
            13'd1417: data <= 8'hFF;
            13'd1418: data <= 8'hFF;
            13'd1419: data <= 8'h80;
            13'd1420: data <= 8'h07;
            13'd1421: data <= 8'hFF;
            13'd1422: data <= 8'hFF;
            13'd1423: data <= 8'hFF;
            13'd1424: data <= 8'hFF;
            13'd1425: data <= 8'hFF;
            13'd1426: data <= 8'hFF;
            13'd1427: data <= 8'hE0;
            13'd1428: data <= 8'h00;
            13'd1429: data <= 8'h00;
            13'd1430: data <= 8'h7F;
            13'd1431: data <= 8'hFF;
            13'd1432: data <= 8'hFF;
            13'd1433: data <= 8'hFF;
            13'd1434: data <= 8'h80;
            13'd1435: data <= 8'h00;
            13'd1436: data <= 8'h00;
            13'd1437: data <= 8'h00;
            13'd1438: data <= 8'h00;
            13'd1439: data <= 8'h00;
            13'd1440: data <= 8'h00;
            13'd1441: data <= 8'h00;
            13'd1442: data <= 8'h00;
            13'd1443: data <= 8'h00;
            13'd1444: data <= 8'h00;
            13'd1445: data <= 8'h03;
            13'd1446: data <= 8'hFF;
            13'd1447: data <= 8'hFF;
            13'd1448: data <= 8'hFF;
            13'd1449: data <= 8'h00;
            13'd1450: data <= 8'h0F;
            13'd1451: data <= 8'hFF;
            13'd1452: data <= 8'hFF;
            13'd1453: data <= 8'hFF;
            13'd1454: data <= 8'hFF;
            13'd1455: data <= 8'hFF;
            13'd1456: data <= 8'hFF;
            13'd1457: data <= 8'hFE;
            13'd1458: data <= 8'h00;
            13'd1459: data <= 8'h00;
            13'd1460: data <= 8'h3F;
            13'd1461: data <= 8'hFF;
            13'd1462: data <= 8'hFF;
            13'd1463: data <= 8'hFF;
            13'd1464: data <= 8'h80;
            13'd1465: data <= 8'h00;
            13'd1466: data <= 8'h00;
            13'd1467: data <= 8'h00;
            13'd1468: data <= 8'h00;
            13'd1469: data <= 8'h00;
            13'd1470: data <= 8'h00;
            13'd1471: data <= 8'h00;
            13'd1472: data <= 8'h00;
            13'd1473: data <= 8'h00;
            13'd1474: data <= 8'h00;
            13'd1475: data <= 8'h03;
            13'd1476: data <= 8'hFF;
            13'd1477: data <= 8'hFF;
            13'd1478: data <= 8'hFE;
            13'd1479: data <= 8'h00;
            13'd1480: data <= 8'h3F;
            13'd1481: data <= 8'hFF;
            13'd1482: data <= 8'hFF;
            13'd1483: data <= 8'hFF;
            13'd1484: data <= 8'hFF;
            13'd1485: data <= 8'hFF;
            13'd1486: data <= 8'hFF;
            13'd1487: data <= 8'hFF;
            13'd1488: data <= 8'h80;
            13'd1489: data <= 8'h00;
            13'd1490: data <= 8'h3F;
            13'd1491: data <= 8'hFF;
            13'd1492: data <= 8'hFF;
            13'd1493: data <= 8'hFF;
            13'd1494: data <= 8'h80;
            13'd1495: data <= 8'h00;
            13'd1496: data <= 8'h00;
            13'd1497: data <= 8'h00;
            13'd1498: data <= 8'h00;
            13'd1499: data <= 8'h00;
            13'd1500: data <= 8'h00;
            13'd1501: data <= 8'h00;
            13'd1502: data <= 8'h00;
            13'd1503: data <= 8'h00;
            13'd1504: data <= 8'h00;
            13'd1505: data <= 8'h03;
            13'd1506: data <= 8'hFF;
            13'd1507: data <= 8'hFF;
            13'd1508: data <= 8'hFC;
            13'd1509: data <= 8'h00;
            13'd1510: data <= 8'hFF;
            13'd1511: data <= 8'hFF;
            13'd1512: data <= 8'hFF;
            13'd1513: data <= 8'hFF;
            13'd1514: data <= 8'hFF;
            13'd1515: data <= 8'hFF;
            13'd1516: data <= 8'hFF;
            13'd1517: data <= 8'hFF;
            13'd1518: data <= 8'hFF;
            13'd1519: data <= 8'hE0;
            13'd1520: data <= 8'h3F;
            13'd1521: data <= 8'hFF;
            13'd1522: data <= 8'hFF;
            13'd1523: data <= 8'hFF;
            13'd1524: data <= 8'h80;
            13'd1525: data <= 8'h00;
            13'd1526: data <= 8'h00;
            13'd1527: data <= 8'h00;
            13'd1528: data <= 8'h00;
            13'd1529: data <= 8'h00;
            13'd1530: data <= 8'h00;
            13'd1531: data <= 8'h00;
            13'd1532: data <= 8'h00;
            13'd1533: data <= 8'h00;
            13'd1534: data <= 8'h00;
            13'd1535: data <= 8'h03;
            13'd1536: data <= 8'hFF;
            13'd1537: data <= 8'hFF;
            13'd1538: data <= 8'hF8;
            13'd1539: data <= 8'h01;
            13'd1540: data <= 8'hFF;
            13'd1541: data <= 8'hFF;
            13'd1542: data <= 8'hFF;
            13'd1543: data <= 8'hFF;
            13'd1544: data <= 8'hFF;
            13'd1545: data <= 8'hFF;
            13'd1546: data <= 8'hFF;
            13'd1547: data <= 8'hFF;
            13'd1548: data <= 8'hFF;
            13'd1549: data <= 8'hF0;
            13'd1550: data <= 8'h1F;
            13'd1551: data <= 8'hFF;
            13'd1552: data <= 8'hFF;
            13'd1553: data <= 8'hFF;
            13'd1554: data <= 8'h80;
            13'd1555: data <= 8'h00;
            13'd1556: data <= 8'h00;
            13'd1557: data <= 8'h00;
            13'd1558: data <= 8'h00;
            13'd1559: data <= 8'h00;
            13'd1560: data <= 8'h00;
            13'd1561: data <= 8'h00;
            13'd1562: data <= 8'h00;
            13'd1563: data <= 8'h00;
            13'd1564: data <= 8'h00;
            13'd1565: data <= 8'h03;
            13'd1566: data <= 8'hFF;
            13'd1567: data <= 8'hFF;
            13'd1568: data <= 8'hF0;
            13'd1569: data <= 8'h03;
            13'd1570: data <= 8'hFF;
            13'd1571: data <= 8'hFF;
            13'd1572: data <= 8'hFF;
            13'd1573: data <= 8'hFF;
            13'd1574: data <= 8'hFF;
            13'd1575: data <= 8'hFF;
            13'd1576: data <= 8'hFF;
            13'd1577: data <= 8'hFF;
            13'd1578: data <= 8'hFF;
            13'd1579: data <= 8'hF0;
            13'd1580: data <= 8'h1F;
            13'd1581: data <= 8'hFF;
            13'd1582: data <= 8'hFF;
            13'd1583: data <= 8'hFF;
            13'd1584: data <= 8'h80;
            13'd1585: data <= 8'h00;
            13'd1586: data <= 8'h00;
            13'd1587: data <= 8'h00;
            13'd1588: data <= 8'h00;
            13'd1589: data <= 8'h00;
            13'd1590: data <= 8'h00;
            13'd1591: data <= 8'h00;
            13'd1592: data <= 8'h00;
            13'd1593: data <= 8'h00;
            13'd1594: data <= 8'h00;
            13'd1595: data <= 8'h03;
            13'd1596: data <= 8'hFF;
            13'd1597: data <= 8'hFF;
            13'd1598: data <= 8'hF0;
            13'd1599: data <= 8'h0F;
            13'd1600: data <= 8'hFF;
            13'd1601: data <= 8'hFF;
            13'd1602: data <= 8'hFF;
            13'd1603: data <= 8'hFF;
            13'd1604: data <= 8'hFF;
            13'd1605: data <= 8'hFF;
            13'd1606: data <= 8'hFF;
            13'd1607: data <= 8'hFF;
            13'd1608: data <= 8'hFF;
            13'd1609: data <= 8'hF0;
            13'd1610: data <= 8'h1F;
            13'd1611: data <= 8'hFF;
            13'd1612: data <= 8'hFF;
            13'd1613: data <= 8'hFF;
            13'd1614: data <= 8'h80;
            13'd1615: data <= 8'h00;
            13'd1616: data <= 8'h00;
            13'd1617: data <= 8'h00;
            13'd1618: data <= 8'h00;
            13'd1619: data <= 8'h00;
            13'd1620: data <= 8'h00;
            13'd1621: data <= 8'h00;
            13'd1622: data <= 8'h00;
            13'd1623: data <= 8'h00;
            13'd1624: data <= 8'h00;
            13'd1625: data <= 8'h03;
            13'd1626: data <= 8'hFF;
            13'd1627: data <= 8'hFF;
            13'd1628: data <= 8'hE0;
            13'd1629: data <= 8'h0F;
            13'd1630: data <= 8'hFF;
            13'd1631: data <= 8'hFF;
            13'd1632: data <= 8'hFF;
            13'd1633: data <= 8'hFF;
            13'd1634: data <= 8'hFF;
            13'd1635: data <= 8'hFF;
            13'd1636: data <= 8'hFF;
            13'd1637: data <= 8'hFF;
            13'd1638: data <= 8'hFF;
            13'd1639: data <= 8'hF8;
            13'd1640: data <= 8'h0F;
            13'd1641: data <= 8'hFF;
            13'd1642: data <= 8'hFF;
            13'd1643: data <= 8'hFF;
            13'd1644: data <= 8'h80;
            13'd1645: data <= 8'h00;
            13'd1646: data <= 8'h00;
            13'd1647: data <= 8'h00;
            13'd1648: data <= 8'h00;
            13'd1649: data <= 8'h00;
            13'd1650: data <= 8'h00;
            13'd1651: data <= 8'h00;
            13'd1652: data <= 8'h00;
            13'd1653: data <= 8'h00;
            13'd1654: data <= 8'h00;
            13'd1655: data <= 8'h03;
            13'd1656: data <= 8'hFF;
            13'd1657: data <= 8'hFF;
            13'd1658: data <= 8'hC0;
            13'd1659: data <= 8'h1F;
            13'd1660: data <= 8'hFF;
            13'd1661: data <= 8'hFF;
            13'd1662: data <= 8'hFF;
            13'd1663: data <= 8'hFF;
            13'd1664: data <= 8'hFF;
            13'd1665: data <= 8'hFF;
            13'd1666: data <= 8'hFF;
            13'd1667: data <= 8'hFF;
            13'd1668: data <= 8'hFF;
            13'd1669: data <= 8'hF8;
            13'd1670: data <= 8'h0F;
            13'd1671: data <= 8'hFF;
            13'd1672: data <= 8'hFF;
            13'd1673: data <= 8'hFF;
            13'd1674: data <= 8'h80;
            13'd1675: data <= 8'h00;
            13'd1676: data <= 8'h00;
            13'd1677: data <= 8'h00;
            13'd1678: data <= 8'h00;
            13'd1679: data <= 8'h00;
            13'd1680: data <= 8'h00;
            13'd1681: data <= 8'h00;
            13'd1682: data <= 8'h00;
            13'd1683: data <= 8'h00;
            13'd1684: data <= 8'h00;
            13'd1685: data <= 8'h03;
            13'd1686: data <= 8'hFF;
            13'd1687: data <= 8'hFF;
            13'd1688: data <= 8'hC0;
            13'd1689: data <= 8'h7F;
            13'd1690: data <= 8'hFF;
            13'd1691: data <= 8'hFF;
            13'd1692: data <= 8'hFF;
            13'd1693: data <= 8'hFF;
            13'd1694: data <= 8'hFF;
            13'd1695: data <= 8'hFF;
            13'd1696: data <= 8'hFF;
            13'd1697: data <= 8'hFF;
            13'd1698: data <= 8'hFF;
            13'd1699: data <= 8'hF8;
            13'd1700: data <= 8'h0F;
            13'd1701: data <= 8'hFF;
            13'd1702: data <= 8'hFF;
            13'd1703: data <= 8'hFF;
            13'd1704: data <= 8'h80;
            13'd1705: data <= 8'h00;
            13'd1706: data <= 8'h00;
            13'd1707: data <= 8'h00;
            13'd1708: data <= 8'h00;
            13'd1709: data <= 8'h00;
            13'd1710: data <= 8'h00;
            13'd1711: data <= 8'h00;
            13'd1712: data <= 8'h00;
            13'd1713: data <= 8'h00;
            13'd1714: data <= 8'h00;
            13'd1715: data <= 8'h03;
            13'd1716: data <= 8'hFF;
            13'd1717: data <= 8'hFF;
            13'd1718: data <= 8'h80;
            13'd1719: data <= 8'h7F;
            13'd1720: data <= 8'hFF;
            13'd1721: data <= 8'hFF;
            13'd1722: data <= 8'hFF;
            13'd1723: data <= 8'hFF;
            13'd1724: data <= 8'hFF;
            13'd1725: data <= 8'hFF;
            13'd1726: data <= 8'hFF;
            13'd1727: data <= 8'hFF;
            13'd1728: data <= 8'hFF;
            13'd1729: data <= 8'hF8;
            13'd1730: data <= 8'h07;
            13'd1731: data <= 8'hFF;
            13'd1732: data <= 8'hFF;
            13'd1733: data <= 8'hFF;
            13'd1734: data <= 8'h80;
            13'd1735: data <= 8'h00;
            13'd1736: data <= 8'h00;
            13'd1737: data <= 8'h00;
            13'd1738: data <= 8'h00;
            13'd1739: data <= 8'h00;
            13'd1740: data <= 8'h00;
            13'd1741: data <= 8'h00;
            13'd1742: data <= 8'h00;
            13'd1743: data <= 8'h00;
            13'd1744: data <= 8'h00;
            13'd1745: data <= 8'h03;
            13'd1746: data <= 8'hFF;
            13'd1747: data <= 8'hFF;
            13'd1748: data <= 8'h80;
            13'd1749: data <= 8'hFF;
            13'd1750: data <= 8'hFF;
            13'd1751: data <= 8'hFF;
            13'd1752: data <= 8'hFF;
            13'd1753: data <= 8'hFF;
            13'd1754: data <= 8'hFF;
            13'd1755: data <= 8'hFF;
            13'd1756: data <= 8'hFF;
            13'd1757: data <= 8'hFF;
            13'd1758: data <= 8'hFF;
            13'd1759: data <= 8'hFC;
            13'd1760: data <= 8'h07;
            13'd1761: data <= 8'hFF;
            13'd1762: data <= 8'hFF;
            13'd1763: data <= 8'hFF;
            13'd1764: data <= 8'h80;
            13'd1765: data <= 8'h00;
            13'd1766: data <= 8'h00;
            13'd1767: data <= 8'h00;
            13'd1768: data <= 8'h00;
            13'd1769: data <= 8'h00;
            13'd1770: data <= 8'h00;
            13'd1771: data <= 8'h00;
            13'd1772: data <= 8'h00;
            13'd1773: data <= 8'h00;
            13'd1774: data <= 8'h00;
            13'd1775: data <= 8'h03;
            13'd1776: data <= 8'hFF;
            13'd1777: data <= 8'hFF;
            13'd1778: data <= 8'h00;
            13'd1779: data <= 8'hFF;
            13'd1780: data <= 8'hFF;
            13'd1781: data <= 8'hFF;
            13'd1782: data <= 8'hFF;
            13'd1783: data <= 8'hFF;
            13'd1784: data <= 8'hFF;
            13'd1785: data <= 8'hFF;
            13'd1786: data <= 8'hFF;
            13'd1787: data <= 8'hFF;
            13'd1788: data <= 8'hFF;
            13'd1789: data <= 8'hFC;
            13'd1790: data <= 8'h07;
            13'd1791: data <= 8'hFF;
            13'd1792: data <= 8'hFF;
            13'd1793: data <= 8'hFF;
            13'd1794: data <= 8'h80;
            13'd1795: data <= 8'h00;
            13'd1796: data <= 8'h00;
            13'd1797: data <= 8'h00;
            13'd1798: data <= 8'h00;
            13'd1799: data <= 8'h00;
            13'd1800: data <= 8'h00;
            13'd1801: data <= 8'h00;
            13'd1802: data <= 8'h00;
            13'd1803: data <= 8'h00;
            13'd1804: data <= 8'h00;
            13'd1805: data <= 8'h03;
            13'd1806: data <= 8'hFF;
            13'd1807: data <= 8'hFF;
            13'd1808: data <= 8'h01;
            13'd1809: data <= 8'hFF;
            13'd1810: data <= 8'hFF;
            13'd1811: data <= 8'hFF;
            13'd1812: data <= 8'hFF;
            13'd1813: data <= 8'hFF;
            13'd1814: data <= 8'hFF;
            13'd1815: data <= 8'hFF;
            13'd1816: data <= 8'hFF;
            13'd1817: data <= 8'hFF;
            13'd1818: data <= 8'hFF;
            13'd1819: data <= 8'hFE;
            13'd1820: data <= 8'h03;
            13'd1821: data <= 8'hFF;
            13'd1822: data <= 8'hFF;
            13'd1823: data <= 8'hFF;
            13'd1824: data <= 8'h80;
            13'd1825: data <= 8'h00;
            13'd1826: data <= 8'h00;
            13'd1827: data <= 8'h00;
            13'd1828: data <= 8'h00;
            13'd1829: data <= 8'h00;
            13'd1830: data <= 8'h00;
            13'd1831: data <= 8'h00;
            13'd1832: data <= 8'h00;
            13'd1833: data <= 8'h00;
            13'd1834: data <= 8'h00;
            13'd1835: data <= 8'h03;
            13'd1836: data <= 8'hFF;
            13'd1837: data <= 8'hFF;
            13'd1838: data <= 8'h01;
            13'd1839: data <= 8'hFF;
            13'd1840: data <= 8'hFF;
            13'd1841: data <= 8'hFF;
            13'd1842: data <= 8'hFF;
            13'd1843: data <= 8'hFF;
            13'd1844: data <= 8'hFF;
            13'd1845: data <= 8'hFF;
            13'd1846: data <= 8'hFF;
            13'd1847: data <= 8'hFF;
            13'd1848: data <= 8'hFF;
            13'd1849: data <= 8'hFE;
            13'd1850: data <= 8'h01;
            13'd1851: data <= 8'hFF;
            13'd1852: data <= 8'hFF;
            13'd1853: data <= 8'hFF;
            13'd1854: data <= 8'h80;
            13'd1855: data <= 8'h00;
            13'd1856: data <= 8'h00;
            13'd1857: data <= 8'h00;
            13'd1858: data <= 8'h00;
            13'd1859: data <= 8'h00;
            13'd1860: data <= 8'h00;
            13'd1861: data <= 8'h00;
            13'd1862: data <= 8'h00;
            13'd1863: data <= 8'h00;
            13'd1864: data <= 8'h00;
            13'd1865: data <= 8'h03;
            13'd1866: data <= 8'hFF;
            13'd1867: data <= 8'hFF;
            13'd1868: data <= 8'h01;
            13'd1869: data <= 8'hFF;
            13'd1870: data <= 8'hF9;
            13'd1871: data <= 8'hFF;
            13'd1872: data <= 8'hFF;
            13'd1873: data <= 8'hFF;
            13'd1874: data <= 8'hFF;
            13'd1875: data <= 8'hFF;
            13'd1876: data <= 8'hFF;
            13'd1877: data <= 8'hFF;
            13'd1878: data <= 8'hFF;
            13'd1879: data <= 8'hFE;
            13'd1880: data <= 8'h01;
            13'd1881: data <= 8'hFF;
            13'd1882: data <= 8'hFF;
            13'd1883: data <= 8'hFF;
            13'd1884: data <= 8'h80;
            13'd1885: data <= 8'h00;
            13'd1886: data <= 8'h00;
            13'd1887: data <= 8'h00;
            13'd1888: data <= 8'h00;
            13'd1889: data <= 8'h00;
            13'd1890: data <= 8'h00;
            13'd1891: data <= 8'h00;
            13'd1892: data <= 8'h00;
            13'd1893: data <= 8'h00;
            13'd1894: data <= 8'h00;
            13'd1895: data <= 8'h03;
            13'd1896: data <= 8'hFF;
            13'd1897: data <= 8'hFE;
            13'd1898: data <= 8'h03;
            13'd1899: data <= 8'hFF;
            13'd1900: data <= 8'hF0;
            13'd1901: data <= 8'hFF;
            13'd1902: data <= 8'hFF;
            13'd1903: data <= 8'hFF;
            13'd1904: data <= 8'hFF;
            13'd1905: data <= 8'hFF;
            13'd1906: data <= 8'hFF;
            13'd1907: data <= 8'hFF;
            13'd1908: data <= 8'hFF;
            13'd1909: data <= 8'hFF;
            13'd1910: data <= 8'h00;
            13'd1911: data <= 8'hFF;
            13'd1912: data <= 8'hFF;
            13'd1913: data <= 8'hFF;
            13'd1914: data <= 8'h80;
            13'd1915: data <= 8'h00;
            13'd1916: data <= 8'h00;
            13'd1917: data <= 8'h00;
            13'd1918: data <= 8'h00;
            13'd1919: data <= 8'h00;
            13'd1920: data <= 8'h00;
            13'd1921: data <= 8'h00;
            13'd1922: data <= 8'h00;
            13'd1923: data <= 8'h00;
            13'd1924: data <= 8'h00;
            13'd1925: data <= 8'h03;
            13'd1926: data <= 8'hFF;
            13'd1927: data <= 8'hFE;
            13'd1928: data <= 8'h03;
            13'd1929: data <= 8'hFF;
            13'd1930: data <= 8'hF0;
            13'd1931: data <= 8'hFF;
            13'd1932: data <= 8'hC7;
            13'd1933: data <= 8'hFF;
            13'd1934: data <= 8'hFF;
            13'd1935: data <= 8'hFF;
            13'd1936: data <= 8'hFF;
            13'd1937: data <= 8'hFF;
            13'd1938: data <= 8'hFF;
            13'd1939: data <= 8'hFF;
            13'd1940: data <= 8'h00;
            13'd1941: data <= 8'hFF;
            13'd1942: data <= 8'hFF;
            13'd1943: data <= 8'hFF;
            13'd1944: data <= 8'h80;
            13'd1945: data <= 8'h00;
            13'd1946: data <= 8'h00;
            13'd1947: data <= 8'h00;
            13'd1948: data <= 8'h00;
            13'd1949: data <= 8'h00;
            13'd1950: data <= 8'h00;
            13'd1951: data <= 8'h00;
            13'd1952: data <= 8'h00;
            13'd1953: data <= 8'h00;
            13'd1954: data <= 8'h00;
            13'd1955: data <= 8'h03;
            13'd1956: data <= 8'hFF;
            13'd1957: data <= 8'hFE;
            13'd1958: data <= 8'h07;
            13'd1959: data <= 8'hFF;
            13'd1960: data <= 8'hF0;
            13'd1961: data <= 8'hFF;
            13'd1962: data <= 8'h83;
            13'd1963: data <= 8'hFF;
            13'd1964: data <= 8'hFF;
            13'd1965: data <= 8'hFF;
            13'd1966: data <= 8'hFF;
            13'd1967: data <= 8'hFF;
            13'd1968: data <= 8'hFF;
            13'd1969: data <= 8'hFF;
            13'd1970: data <= 8'h80;
            13'd1971: data <= 8'h7F;
            13'd1972: data <= 8'hFF;
            13'd1973: data <= 8'hFF;
            13'd1974: data <= 8'h80;
            13'd1975: data <= 8'h00;
            13'd1976: data <= 8'h00;
            13'd1977: data <= 8'h00;
            13'd1978: data <= 8'h00;
            13'd1979: data <= 8'h00;
            13'd1980: data <= 8'h00;
            13'd1981: data <= 8'h00;
            13'd1982: data <= 8'h00;
            13'd1983: data <= 8'h00;
            13'd1984: data <= 8'h00;
            13'd1985: data <= 8'h03;
            13'd1986: data <= 8'hFF;
            13'd1987: data <= 8'hFE;
            13'd1988: data <= 8'h07;
            13'd1989: data <= 8'hFF;
            13'd1990: data <= 8'hFD;
            13'd1991: data <= 8'hFF;
            13'd1992: data <= 8'h83;
            13'd1993: data <= 8'hFF;
            13'd1994: data <= 8'hFF;
            13'd1995: data <= 8'hFF;
            13'd1996: data <= 8'hFF;
            13'd1997: data <= 8'hFF;
            13'd1998: data <= 8'hFF;
            13'd1999: data <= 8'hFF;
            13'd2000: data <= 8'h80;
            13'd2001: data <= 8'h7F;
            13'd2002: data <= 8'hFF;
            13'd2003: data <= 8'hFF;
            13'd2004: data <= 8'h80;
            13'd2005: data <= 8'h00;
            13'd2006: data <= 8'h00;
            13'd2007: data <= 8'h00;
            13'd2008: data <= 8'h00;
            13'd2009: data <= 8'h00;
            13'd2010: data <= 8'h00;
            13'd2011: data <= 8'h00;
            13'd2012: data <= 8'h00;
            13'd2013: data <= 8'h00;
            13'd2014: data <= 8'h00;
            13'd2015: data <= 8'h03;
            13'd2016: data <= 8'hFF;
            13'd2017: data <= 8'hFE;
            13'd2018: data <= 8'h07;
            13'd2019: data <= 8'hFF;
            13'd2020: data <= 8'hFF;
            13'd2021: data <= 8'hFF;
            13'd2022: data <= 8'h83;
            13'd2023: data <= 8'hFF;
            13'd2024: data <= 8'hFF;
            13'd2025: data <= 8'hFF;
            13'd2026: data <= 8'hFF;
            13'd2027: data <= 8'hFF;
            13'd2028: data <= 8'hFF;
            13'd2029: data <= 8'hFF;
            13'd2030: data <= 8'hC0;
            13'd2031: data <= 8'h3F;
            13'd2032: data <= 8'hFF;
            13'd2033: data <= 8'hFF;
            13'd2034: data <= 8'h80;
            13'd2035: data <= 8'h00;
            13'd2036: data <= 8'h00;
            13'd2037: data <= 8'h00;
            13'd2038: data <= 8'h00;
            13'd2039: data <= 8'h00;
            13'd2040: data <= 8'h00;
            13'd2041: data <= 8'h00;
            13'd2042: data <= 8'h00;
            13'd2043: data <= 8'h00;
            13'd2044: data <= 8'h00;
            13'd2045: data <= 8'h03;
            13'd2046: data <= 8'hFF;
            13'd2047: data <= 8'hFE;
            13'd2048: data <= 8'h07;
            13'd2049: data <= 8'hFF;
            13'd2050: data <= 8'hFF;
            13'd2051: data <= 8'hFF;
            13'd2052: data <= 8'hEF;
            13'd2053: data <= 8'hFF;
            13'd2054: data <= 8'hFF;
            13'd2055: data <= 8'hFF;
            13'd2056: data <= 8'hFF;
            13'd2057: data <= 8'hFF;
            13'd2058: data <= 8'hFF;
            13'd2059: data <= 8'hFF;
            13'd2060: data <= 8'hE0;
            13'd2061: data <= 8'h3F;
            13'd2062: data <= 8'hFF;
            13'd2063: data <= 8'hFF;
            13'd2064: data <= 8'h80;
            13'd2065: data <= 8'h00;
            13'd2066: data <= 8'h00;
            13'd2067: data <= 8'h00;
            13'd2068: data <= 8'h00;
            13'd2069: data <= 8'h00;
            13'd2070: data <= 8'h00;
            13'd2071: data <= 8'h00;
            13'd2072: data <= 8'h00;
            13'd2073: data <= 8'h00;
            13'd2074: data <= 8'h00;
            13'd2075: data <= 8'h03;
            13'd2076: data <= 8'hFF;
            13'd2077: data <= 8'hFE;
            13'd2078: data <= 8'h07;
            13'd2079: data <= 8'hFF;
            13'd2080: data <= 8'hFF;
            13'd2081: data <= 8'hFF;
            13'd2082: data <= 8'hFF;
            13'd2083: data <= 8'hFF;
            13'd2084: data <= 8'hFF;
            13'd2085: data <= 8'hFF;
            13'd2086: data <= 8'hFF;
            13'd2087: data <= 8'hFF;
            13'd2088: data <= 8'hFF;
            13'd2089: data <= 8'hFF;
            13'd2090: data <= 8'hE0;
            13'd2091: data <= 8'h1F;
            13'd2092: data <= 8'hFF;
            13'd2093: data <= 8'hFF;
            13'd2094: data <= 8'h80;
            13'd2095: data <= 8'h00;
            13'd2096: data <= 8'h00;
            13'd2097: data <= 8'h00;
            13'd2098: data <= 8'h00;
            13'd2099: data <= 8'h00;
            13'd2100: data <= 8'h00;
            13'd2101: data <= 8'h00;
            13'd2102: data <= 8'h00;
            13'd2103: data <= 8'h00;
            13'd2104: data <= 8'h00;
            13'd2105: data <= 8'h03;
            13'd2106: data <= 8'hFF;
            13'd2107: data <= 8'hFE;
            13'd2108: data <= 8'h07;
            13'd2109: data <= 8'hFF;
            13'd2110: data <= 8'hFF;
            13'd2111: data <= 8'hFF;
            13'd2112: data <= 8'hFF;
            13'd2113: data <= 8'hFF;
            13'd2114: data <= 8'hFF;
            13'd2115: data <= 8'hFF;
            13'd2116: data <= 8'hFF;
            13'd2117: data <= 8'hFF;
            13'd2118: data <= 8'hFF;
            13'd2119: data <= 8'hFF;
            13'd2120: data <= 8'hF0;
            13'd2121: data <= 8'h0F;
            13'd2122: data <= 8'hFF;
            13'd2123: data <= 8'hFF;
            13'd2124: data <= 8'h80;
            13'd2125: data <= 8'h00;
            13'd2126: data <= 8'h00;
            13'd2127: data <= 8'h00;
            13'd2128: data <= 8'h00;
            13'd2129: data <= 8'h00;
            13'd2130: data <= 8'h00;
            13'd2131: data <= 8'h00;
            13'd2132: data <= 8'h00;
            13'd2133: data <= 8'h00;
            13'd2134: data <= 8'h00;
            13'd2135: data <= 8'h03;
            13'd2136: data <= 8'hFF;
            13'd2137: data <= 8'hFE;
            13'd2138: data <= 8'h07;
            13'd2139: data <= 8'hFF;
            13'd2140: data <= 8'hFF;
            13'd2141: data <= 8'hFF;
            13'd2142: data <= 8'hFF;
            13'd2143: data <= 8'hFF;
            13'd2144: data <= 8'hFF;
            13'd2145: data <= 8'hFF;
            13'd2146: data <= 8'hFF;
            13'd2147: data <= 8'hFF;
            13'd2148: data <= 8'hFF;
            13'd2149: data <= 8'hFF;
            13'd2150: data <= 8'hF0;
            13'd2151: data <= 8'h0F;
            13'd2152: data <= 8'hFF;
            13'd2153: data <= 8'hFF;
            13'd2154: data <= 8'h80;
            13'd2155: data <= 8'h00;
            13'd2156: data <= 8'h00;
            13'd2157: data <= 8'h00;
            13'd2158: data <= 8'h00;
            13'd2159: data <= 8'h00;
            13'd2160: data <= 8'h00;
            13'd2161: data <= 8'h00;
            13'd2162: data <= 8'h00;
            13'd2163: data <= 8'h00;
            13'd2164: data <= 8'h00;
            13'd2165: data <= 8'h03;
            13'd2166: data <= 8'hFF;
            13'd2167: data <= 8'hFE;
            13'd2168: data <= 8'h07;
            13'd2169: data <= 8'hFF;
            13'd2170: data <= 8'hFF;
            13'd2171: data <= 8'hFF;
            13'd2172: data <= 8'hFF;
            13'd2173: data <= 8'hFF;
            13'd2174: data <= 8'hFF;
            13'd2175: data <= 8'hFF;
            13'd2176: data <= 8'hFF;
            13'd2177: data <= 8'hFF;
            13'd2178: data <= 8'hFF;
            13'd2179: data <= 8'hFF;
            13'd2180: data <= 8'hF8;
            13'd2181: data <= 8'h0F;
            13'd2182: data <= 8'hFF;
            13'd2183: data <= 8'hFF;
            13'd2184: data <= 8'h80;
            13'd2185: data <= 8'h00;
            13'd2186: data <= 8'h00;
            13'd2187: data <= 8'h00;
            13'd2188: data <= 8'h00;
            13'd2189: data <= 8'h00;
            13'd2190: data <= 8'h00;
            13'd2191: data <= 8'h00;
            13'd2192: data <= 8'h00;
            13'd2193: data <= 8'h00;
            13'd2194: data <= 8'h00;
            13'd2195: data <= 8'h03;
            13'd2196: data <= 8'hFF;
            13'd2197: data <= 8'hFE;
            13'd2198: data <= 8'h07;
            13'd2199: data <= 8'hFF;
            13'd2200: data <= 8'hFF;
            13'd2201: data <= 8'hFF;
            13'd2202: data <= 8'hFF;
            13'd2203: data <= 8'hFF;
            13'd2204: data <= 8'hFF;
            13'd2205: data <= 8'hFF;
            13'd2206: data <= 8'hFF;
            13'd2207: data <= 8'hFF;
            13'd2208: data <= 8'hFF;
            13'd2209: data <= 8'hFF;
            13'd2210: data <= 8'hFC;
            13'd2211: data <= 8'h07;
            13'd2212: data <= 8'hFF;
            13'd2213: data <= 8'hFF;
            13'd2214: data <= 8'h80;
            13'd2215: data <= 8'h00;
            13'd2216: data <= 8'h00;
            13'd2217: data <= 8'h00;
            13'd2218: data <= 8'h00;
            13'd2219: data <= 8'h00;
            13'd2220: data <= 8'h00;
            13'd2221: data <= 8'h00;
            13'd2222: data <= 8'h00;
            13'd2223: data <= 8'h00;
            13'd2224: data <= 8'h00;
            13'd2225: data <= 8'h03;
            13'd2226: data <= 8'hFF;
            13'd2227: data <= 8'hFE;
            13'd2228: data <= 8'h07;
            13'd2229: data <= 8'hFF;
            13'd2230: data <= 8'hFB;
            13'd2231: data <= 8'hFF;
            13'd2232: data <= 8'hFF;
            13'd2233: data <= 8'hFF;
            13'd2234: data <= 8'hFF;
            13'd2235: data <= 8'hFF;
            13'd2236: data <= 8'hFF;
            13'd2237: data <= 8'hFF;
            13'd2238: data <= 8'hFF;
            13'd2239: data <= 8'hFF;
            13'd2240: data <= 8'hFC;
            13'd2241: data <= 8'h07;
            13'd2242: data <= 8'hFF;
            13'd2243: data <= 8'hFF;
            13'd2244: data <= 8'h80;
            13'd2245: data <= 8'h00;
            13'd2246: data <= 8'h00;
            13'd2247: data <= 8'h00;
            13'd2248: data <= 8'h00;
            13'd2249: data <= 8'h00;
            13'd2250: data <= 8'h00;
            13'd2251: data <= 8'h00;
            13'd2252: data <= 8'h00;
            13'd2253: data <= 8'h00;
            13'd2254: data <= 8'h00;
            13'd2255: data <= 8'h03;
            13'd2256: data <= 8'hFF;
            13'd2257: data <= 8'hFF;
            13'd2258: data <= 8'h03;
            13'd2259: data <= 8'hFF;
            13'd2260: data <= 8'hF1;
            13'd2261: data <= 8'hFF;
            13'd2262: data <= 8'hFF;
            13'd2263: data <= 8'hFF;
            13'd2264: data <= 8'hFF;
            13'd2265: data <= 8'hFF;
            13'd2266: data <= 8'hFF;
            13'd2267: data <= 8'hFF;
            13'd2268: data <= 8'hFF;
            13'd2269: data <= 8'hFF;
            13'd2270: data <= 8'hFE;
            13'd2271: data <= 8'h03;
            13'd2272: data <= 8'hFF;
            13'd2273: data <= 8'hFF;
            13'd2274: data <= 8'h80;
            13'd2275: data <= 8'h00;
            13'd2276: data <= 8'h00;
            13'd2277: data <= 8'h00;
            13'd2278: data <= 8'h00;
            13'd2279: data <= 8'h00;
            13'd2280: data <= 8'h00;
            13'd2281: data <= 8'h00;
            13'd2282: data <= 8'h00;
            13'd2283: data <= 8'h00;
            13'd2284: data <= 8'h00;
            13'd2285: data <= 8'h03;
            13'd2286: data <= 8'hFF;
            13'd2287: data <= 8'hFF;
            13'd2288: data <= 8'h03;
            13'd2289: data <= 8'hFF;
            13'd2290: data <= 8'hE0;
            13'd2291: data <= 8'h38;
            13'd2292: data <= 8'h3F;
            13'd2293: data <= 8'hFF;
            13'd2294: data <= 8'hFF;
            13'd2295: data <= 8'hFF;
            13'd2296: data <= 8'hFF;
            13'd2297: data <= 8'hFF;
            13'd2298: data <= 8'hFF;
            13'd2299: data <= 8'hFF;
            13'd2300: data <= 8'hFE;
            13'd2301: data <= 8'h03;
            13'd2302: data <= 8'hFF;
            13'd2303: data <= 8'hFF;
            13'd2304: data <= 8'h80;
            13'd2305: data <= 8'h00;
            13'd2306: data <= 8'h00;
            13'd2307: data <= 8'h00;
            13'd2308: data <= 8'h00;
            13'd2309: data <= 8'h00;
            13'd2310: data <= 8'h00;
            13'd2311: data <= 8'h00;
            13'd2312: data <= 8'h00;
            13'd2313: data <= 8'h00;
            13'd2314: data <= 8'h00;
            13'd2315: data <= 8'h03;
            13'd2316: data <= 8'hFF;
            13'd2317: data <= 8'hFF;
            13'd2318: data <= 8'h83;
            13'd2319: data <= 8'hFF;
            13'd2320: data <= 8'hE0;
            13'd2321: data <= 8'h00;
            13'd2322: data <= 8'h3F;
            13'd2323: data <= 8'hFF;
            13'd2324: data <= 8'hFF;
            13'd2325: data <= 8'hFF;
            13'd2326: data <= 8'hFF;
            13'd2327: data <= 8'hFF;
            13'd2328: data <= 8'hFF;
            13'd2329: data <= 8'hFF;
            13'd2330: data <= 8'hFF;
            13'd2331: data <= 8'h01;
            13'd2332: data <= 8'hFF;
            13'd2333: data <= 8'hFF;
            13'd2334: data <= 8'h80;
            13'd2335: data <= 8'h00;
            13'd2336: data <= 8'h00;
            13'd2337: data <= 8'h00;
            13'd2338: data <= 8'h00;
            13'd2339: data <= 8'h00;
            13'd2340: data <= 8'h00;
            13'd2341: data <= 8'h00;
            13'd2342: data <= 8'h00;
            13'd2343: data <= 8'h00;
            13'd2344: data <= 8'h00;
            13'd2345: data <= 8'h03;
            13'd2346: data <= 8'hFF;
            13'd2347: data <= 8'hFF;
            13'd2348: data <= 8'h81;
            13'd2349: data <= 8'h03;
            13'd2350: data <= 8'hE0;
            13'd2351: data <= 8'h00;
            13'd2352: data <= 8'h3F;
            13'd2353: data <= 8'hFF;
            13'd2354: data <= 8'hFF;
            13'd2355: data <= 8'hFF;
            13'd2356: data <= 8'hFF;
            13'd2357: data <= 8'hFF;
            13'd2358: data <= 8'hFF;
            13'd2359: data <= 8'hFF;
            13'd2360: data <= 8'hFF;
            13'd2361: data <= 8'h00;
            13'd2362: data <= 8'hFF;
            13'd2363: data <= 8'hFF;
            13'd2364: data <= 8'h80;
            13'd2365: data <= 8'h00;
            13'd2366: data <= 8'h00;
            13'd2367: data <= 8'h00;
            13'd2368: data <= 8'h00;
            13'd2369: data <= 8'h00;
            13'd2370: data <= 8'h00;
            13'd2371: data <= 8'h00;
            13'd2372: data <= 8'h00;
            13'd2373: data <= 8'h00;
            13'd2374: data <= 8'h00;
            13'd2375: data <= 8'h03;
            13'd2376: data <= 8'hFF;
            13'd2377: data <= 8'hFF;
            13'd2378: data <= 8'hC0;
            13'd2379: data <= 8'h00;
            13'd2380: data <= 8'h70;
            13'd2381: data <= 8'h00;
            13'd2382: data <= 8'h1F;
            13'd2383: data <= 8'hFF;
            13'd2384: data <= 8'hFF;
            13'd2385: data <= 8'hFF;
            13'd2386: data <= 8'hFF;
            13'd2387: data <= 8'hFF;
            13'd2388: data <= 8'hFF;
            13'd2389: data <= 8'hFF;
            13'd2390: data <= 8'hFF;
            13'd2391: data <= 8'h80;
            13'd2392: data <= 8'h7F;
            13'd2393: data <= 8'hFF;
            13'd2394: data <= 8'h80;
            13'd2395: data <= 8'h00;
            13'd2396: data <= 8'h00;
            13'd2397: data <= 8'h00;
            13'd2398: data <= 8'h00;
            13'd2399: data <= 8'h00;
            13'd2400: data <= 8'h00;
            13'd2401: data <= 8'h00;
            13'd2402: data <= 8'h00;
            13'd2403: data <= 8'h00;
            13'd2404: data <= 8'h00;
            13'd2405: data <= 8'h03;
            13'd2406: data <= 8'hFF;
            13'd2407: data <= 8'hFF;
            13'd2408: data <= 8'hE0;
            13'd2409: data <= 8'h00;
            13'd2410: data <= 8'h18;
            13'd2411: data <= 8'h00;
            13'd2412: data <= 8'h7F;
            13'd2413: data <= 8'hFF;
            13'd2414: data <= 8'hFF;
            13'd2415: data <= 8'hFF;
            13'd2416: data <= 8'hFF;
            13'd2417: data <= 8'hFF;
            13'd2418: data <= 8'hFF;
            13'd2419: data <= 8'hFF;
            13'd2420: data <= 8'hFF;
            13'd2421: data <= 8'h80;
            13'd2422: data <= 8'h7F;
            13'd2423: data <= 8'hFF;
            13'd2424: data <= 8'h80;
            13'd2425: data <= 8'h00;
            13'd2426: data <= 8'h00;
            13'd2427: data <= 8'h00;
            13'd2428: data <= 8'h00;
            13'd2429: data <= 8'h00;
            13'd2430: data <= 8'h00;
            13'd2431: data <= 8'h00;
            13'd2432: data <= 8'h00;
            13'd2433: data <= 8'h00;
            13'd2434: data <= 8'h00;
            13'd2435: data <= 8'h03;
            13'd2436: data <= 8'hFF;
            13'd2437: data <= 8'hFF;
            13'd2438: data <= 8'hC0;
            13'd2439: data <= 8'h00;
            13'd2440: data <= 8'h03;
            13'd2441: data <= 8'hF3;
            13'd2442: data <= 8'hFF;
            13'd2443: data <= 8'hFF;
            13'd2444: data <= 8'hFF;
            13'd2445: data <= 8'hFF;
            13'd2446: data <= 8'hFF;
            13'd2447: data <= 8'hFF;
            13'd2448: data <= 8'hFF;
            13'd2449: data <= 8'hFF;
            13'd2450: data <= 8'hFF;
            13'd2451: data <= 8'hC0;
            13'd2452: data <= 8'h7F;
            13'd2453: data <= 8'hFF;
            13'd2454: data <= 8'h80;
            13'd2455: data <= 8'h00;
            13'd2456: data <= 8'h00;
            13'd2457: data <= 8'h00;
            13'd2458: data <= 8'h00;
            13'd2459: data <= 8'h00;
            13'd2460: data <= 8'h00;
            13'd2461: data <= 8'h00;
            13'd2462: data <= 8'h00;
            13'd2463: data <= 8'h00;
            13'd2464: data <= 8'h00;
            13'd2465: data <= 8'h03;
            13'd2466: data <= 8'hFF;
            13'd2467: data <= 8'hFF;
            13'd2468: data <= 8'hC0;
            13'd2469: data <= 8'h00;
            13'd2470: data <= 8'h01;
            13'd2471: data <= 8'hFF;
            13'd2472: data <= 8'hF8;
            13'd2473: data <= 8'h7F;
            13'd2474: data <= 8'hFF;
            13'd2475: data <= 8'hFF;
            13'd2476: data <= 8'hFF;
            13'd2477: data <= 8'hFF;
            13'd2478: data <= 8'hFF;
            13'd2479: data <= 8'hFF;
            13'd2480: data <= 8'hFF;
            13'd2481: data <= 8'hC0;
            13'd2482: data <= 8'h3F;
            13'd2483: data <= 8'hFF;
            13'd2484: data <= 8'h80;
            13'd2485: data <= 8'h00;
            13'd2486: data <= 8'h00;
            13'd2487: data <= 8'h00;
            13'd2488: data <= 8'h00;
            13'd2489: data <= 8'h00;
            13'd2490: data <= 8'h00;
            13'd2491: data <= 8'h00;
            13'd2492: data <= 8'h00;
            13'd2493: data <= 8'h00;
            13'd2494: data <= 8'h00;
            13'd2495: data <= 8'h03;
            13'd2496: data <= 8'hFF;
            13'd2497: data <= 8'hFF;
            13'd2498: data <= 8'hF0;
            13'd2499: data <= 8'h00;
            13'd2500: data <= 8'h00;
            13'd2501: data <= 8'h0F;
            13'd2502: data <= 8'hC0;
            13'd2503: data <= 8'h7F;
            13'd2504: data <= 8'hFF;
            13'd2505: data <= 8'hFF;
            13'd2506: data <= 8'hFF;
            13'd2507: data <= 8'hFF;
            13'd2508: data <= 8'hFF;
            13'd2509: data <= 8'hFF;
            13'd2510: data <= 8'hFF;
            13'd2511: data <= 8'hE0;
            13'd2512: data <= 8'h3F;
            13'd2513: data <= 8'hFF;
            13'd2514: data <= 8'h80;
            13'd2515: data <= 8'h00;
            13'd2516: data <= 8'h00;
            13'd2517: data <= 8'h00;
            13'd2518: data <= 8'h00;
            13'd2519: data <= 8'h00;
            13'd2520: data <= 8'h00;
            13'd2521: data <= 8'h00;
            13'd2522: data <= 8'h00;
            13'd2523: data <= 8'h00;
            13'd2524: data <= 8'h00;
            13'd2525: data <= 8'h03;
            13'd2526: data <= 8'hFF;
            13'd2527: data <= 8'hFF;
            13'd2528: data <= 8'hF8;
            13'd2529: data <= 8'h00;
            13'd2530: data <= 8'h00;
            13'd2531: data <= 8'h04;
            13'd2532: data <= 8'h00;
            13'd2533: data <= 8'h7F;
            13'd2534: data <= 8'hFF;
            13'd2535: data <= 8'hFF;
            13'd2536: data <= 8'hFF;
            13'd2537: data <= 8'hFF;
            13'd2538: data <= 8'hFF;
            13'd2539: data <= 8'hFF;
            13'd2540: data <= 8'hFF;
            13'd2541: data <= 8'hE0;
            13'd2542: data <= 8'h1F;
            13'd2543: data <= 8'hFF;
            13'd2544: data <= 8'h80;
            13'd2545: data <= 8'h00;
            13'd2546: data <= 8'h00;
            13'd2547: data <= 8'h00;
            13'd2548: data <= 8'h00;
            13'd2549: data <= 8'h00;
            13'd2550: data <= 8'h00;
            13'd2551: data <= 8'h00;
            13'd2552: data <= 8'h00;
            13'd2553: data <= 8'h00;
            13'd2554: data <= 8'h00;
            13'd2555: data <= 8'h03;
            13'd2556: data <= 8'hFF;
            13'd2557: data <= 8'hFF;
            13'd2558: data <= 8'hF8;
            13'd2559: data <= 8'h00;
            13'd2560: data <= 8'h00;
            13'd2561: data <= 8'h00;
            13'd2562: data <= 8'h00;
            13'd2563: data <= 8'hFF;
            13'd2564: data <= 8'hFF;
            13'd2565: data <= 8'hFF;
            13'd2566: data <= 8'hFF;
            13'd2567: data <= 8'hFF;
            13'd2568: data <= 8'hFF;
            13'd2569: data <= 8'hFF;
            13'd2570: data <= 8'hFF;
            13'd2571: data <= 8'hF0;
            13'd2572: data <= 8'h1F;
            13'd2573: data <= 8'hFF;
            13'd2574: data <= 8'h80;
            13'd2575: data <= 8'h00;
            13'd2576: data <= 8'h00;
            13'd2577: data <= 8'h00;
            13'd2578: data <= 8'h00;
            13'd2579: data <= 8'h00;
            13'd2580: data <= 8'h00;
            13'd2581: data <= 8'h00;
            13'd2582: data <= 8'h00;
            13'd2583: data <= 8'h00;
            13'd2584: data <= 8'h00;
            13'd2585: data <= 8'h03;
            13'd2586: data <= 8'hFF;
            13'd2587: data <= 8'hFF;
            13'd2588: data <= 8'hFE;
            13'd2589: data <= 8'h00;
            13'd2590: data <= 8'h08;
            13'd2591: data <= 8'h00;
            13'd2592: data <= 8'h01;
            13'd2593: data <= 8'hFF;
            13'd2594: data <= 8'hFF;
            13'd2595: data <= 8'hFF;
            13'd2596: data <= 8'hFF;
            13'd2597: data <= 8'hFF;
            13'd2598: data <= 8'hFF;
            13'd2599: data <= 8'hFF;
            13'd2600: data <= 8'hFF;
            13'd2601: data <= 8'hF0;
            13'd2602: data <= 8'h1F;
            13'd2603: data <= 8'hFF;
            13'd2604: data <= 8'h80;
            13'd2605: data <= 8'h00;
            13'd2606: data <= 8'h00;
            13'd2607: data <= 8'h00;
            13'd2608: data <= 8'h00;
            13'd2609: data <= 8'h00;
            13'd2610: data <= 8'h00;
            13'd2611: data <= 8'h00;
            13'd2612: data <= 8'h00;
            13'd2613: data <= 8'h00;
            13'd2614: data <= 8'h00;
            13'd2615: data <= 8'h03;
            13'd2616: data <= 8'hFF;
            13'd2617: data <= 8'hFF;
            13'd2618: data <= 8'hFF;
            13'd2619: data <= 8'h00;
            13'd2620: data <= 8'h04;
            13'd2621: data <= 8'h00;
            13'd2622: data <= 8'h01;
            13'd2623: data <= 8'hFF;
            13'd2624: data <= 8'hFF;
            13'd2625: data <= 8'hFF;
            13'd2626: data <= 8'hFF;
            13'd2627: data <= 8'hFF;
            13'd2628: data <= 8'hFF;
            13'd2629: data <= 8'hFF;
            13'd2630: data <= 8'hFF;
            13'd2631: data <= 8'hF8;
            13'd2632: data <= 8'h0F;
            13'd2633: data <= 8'hFF;
            13'd2634: data <= 8'h80;
            13'd2635: data <= 8'h00;
            13'd2636: data <= 8'h00;
            13'd2637: data <= 8'h00;
            13'd2638: data <= 8'h00;
            13'd2639: data <= 8'h00;
            13'd2640: data <= 8'h00;
            13'd2641: data <= 8'h00;
            13'd2642: data <= 8'h00;
            13'd2643: data <= 8'h00;
            13'd2644: data <= 8'h00;
            13'd2645: data <= 8'h03;
            13'd2646: data <= 8'hFF;
            13'd2647: data <= 8'hFF;
            13'd2648: data <= 8'hFF;
            13'd2649: data <= 8'h80;
            13'd2650: data <= 8'h07;
            13'd2651: data <= 8'h80;
            13'd2652: data <= 8'h03;
            13'd2653: data <= 8'hFF;
            13'd2654: data <= 8'hFF;
            13'd2655: data <= 8'hFF;
            13'd2656: data <= 8'hFF;
            13'd2657: data <= 8'hFF;
            13'd2658: data <= 8'hFF;
            13'd2659: data <= 8'hFF;
            13'd2660: data <= 8'hFF;
            13'd2661: data <= 8'hF8;
            13'd2662: data <= 8'h0F;
            13'd2663: data <= 8'hFF;
            13'd2664: data <= 8'h80;
            13'd2665: data <= 8'h00;
            13'd2666: data <= 8'h00;
            13'd2667: data <= 8'h00;
            13'd2668: data <= 8'h00;
            13'd2669: data <= 8'h00;
            13'd2670: data <= 8'h00;
            13'd2671: data <= 8'h00;
            13'd2672: data <= 8'h00;
            13'd2673: data <= 8'h00;
            13'd2674: data <= 8'h00;
            13'd2675: data <= 8'h03;
            13'd2676: data <= 8'hFF;
            13'd2677: data <= 8'hFF;
            13'd2678: data <= 8'hFF;
            13'd2679: data <= 8'hE0;
            13'd2680: data <= 8'h07;
            13'd2681: data <= 8'hFF;
            13'd2682: data <= 8'hC7;
            13'd2683: data <= 8'hFF;
            13'd2684: data <= 8'hFF;
            13'd2685: data <= 8'hFF;
            13'd2686: data <= 8'hFF;
            13'd2687: data <= 8'hFF;
            13'd2688: data <= 8'hFF;
            13'd2689: data <= 8'hFF;
            13'd2690: data <= 8'hFF;
            13'd2691: data <= 8'hFC;
            13'd2692: data <= 8'h07;
            13'd2693: data <= 8'hFF;
            13'd2694: data <= 8'h80;
            13'd2695: data <= 8'h00;
            13'd2696: data <= 8'h00;
            13'd2697: data <= 8'h00;
            13'd2698: data <= 8'h00;
            13'd2699: data <= 8'h00;
            13'd2700: data <= 8'h00;
            13'd2701: data <= 8'h00;
            13'd2702: data <= 8'h00;
            13'd2703: data <= 8'h00;
            13'd2704: data <= 8'h00;
            13'd2705: data <= 8'h03;
            13'd2706: data <= 8'hFF;
            13'd2707: data <= 8'hFF;
            13'd2708: data <= 8'hFF;
            13'd2709: data <= 8'hF0;
            13'd2710: data <= 8'h83;
            13'd2711: data <= 8'hFF;
            13'd2712: data <= 8'hC7;
            13'd2713: data <= 8'hFF;
            13'd2714: data <= 8'hFF;
            13'd2715: data <= 8'hFF;
            13'd2716: data <= 8'hFF;
            13'd2717: data <= 8'hFF;
            13'd2718: data <= 8'hFF;
            13'd2719: data <= 8'hFF;
            13'd2720: data <= 8'hFF;
            13'd2721: data <= 8'hFC;
            13'd2722: data <= 8'h07;
            13'd2723: data <= 8'hFF;
            13'd2724: data <= 8'h80;
            13'd2725: data <= 8'h00;
            13'd2726: data <= 8'h00;
            13'd2727: data <= 8'h00;
            13'd2728: data <= 8'h00;
            13'd2729: data <= 8'h00;
            13'd2730: data <= 8'h00;
            13'd2731: data <= 8'h00;
            13'd2732: data <= 8'h00;
            13'd2733: data <= 8'h00;
            13'd2734: data <= 8'h00;
            13'd2735: data <= 8'h03;
            13'd2736: data <= 8'hFF;
            13'd2737: data <= 8'hFF;
            13'd2738: data <= 8'hFF;
            13'd2739: data <= 8'hF0;
            13'd2740: data <= 8'hC1;
            13'd2741: data <= 8'hFF;
            13'd2742: data <= 8'hC7;
            13'd2743: data <= 8'hFF;
            13'd2744: data <= 8'hFF;
            13'd2745: data <= 8'hFF;
            13'd2746: data <= 8'hFF;
            13'd2747: data <= 8'hFF;
            13'd2748: data <= 8'hFF;
            13'd2749: data <= 8'hFF;
            13'd2750: data <= 8'hFF;
            13'd2751: data <= 8'hFC;
            13'd2752: data <= 8'h07;
            13'd2753: data <= 8'hFF;
            13'd2754: data <= 8'h80;
            13'd2755: data <= 8'h00;
            13'd2756: data <= 8'h00;
            13'd2757: data <= 8'h00;
            13'd2758: data <= 8'h00;
            13'd2759: data <= 8'h00;
            13'd2760: data <= 8'h00;
            13'd2761: data <= 8'h00;
            13'd2762: data <= 8'h00;
            13'd2763: data <= 8'h00;
            13'd2764: data <= 8'h00;
            13'd2765: data <= 8'h03;
            13'd2766: data <= 8'hFF;
            13'd2767: data <= 8'hFF;
            13'd2768: data <= 8'hFF;
            13'd2769: data <= 8'hF0;
            13'd2770: data <= 8'hE1;
            13'd2771: data <= 8'hFF;
            13'd2772: data <= 8'hC7;
            13'd2773: data <= 8'hFF;
            13'd2774: data <= 8'hFF;
            13'd2775: data <= 8'hFF;
            13'd2776: data <= 8'hFF;
            13'd2777: data <= 8'hFF;
            13'd2778: data <= 8'hFF;
            13'd2779: data <= 8'hFF;
            13'd2780: data <= 8'hFF;
            13'd2781: data <= 8'hFE;
            13'd2782: data <= 8'h03;
            13'd2783: data <= 8'hFF;
            13'd2784: data <= 8'h80;
            13'd2785: data <= 8'h00;
            13'd2786: data <= 8'h00;
            13'd2787: data <= 8'h00;
            13'd2788: data <= 8'h00;
            13'd2789: data <= 8'h00;
            13'd2790: data <= 8'h00;
            13'd2791: data <= 8'h00;
            13'd2792: data <= 8'h00;
            13'd2793: data <= 8'h00;
            13'd2794: data <= 8'h00;
            13'd2795: data <= 8'h03;
            13'd2796: data <= 8'hFF;
            13'd2797: data <= 8'hFF;
            13'd2798: data <= 8'hFF;
            13'd2799: data <= 8'hF0;
            13'd2800: data <= 8'hF0;
            13'd2801: data <= 8'hFF;
            13'd2802: data <= 8'hC7;
            13'd2803: data <= 8'hFF;
            13'd2804: data <= 8'hFF;
            13'd2805: data <= 8'hFF;
            13'd2806: data <= 8'hFF;
            13'd2807: data <= 8'hFF;
            13'd2808: data <= 8'hFF;
            13'd2809: data <= 8'hFF;
            13'd2810: data <= 8'hFF;
            13'd2811: data <= 8'hFE;
            13'd2812: data <= 8'h03;
            13'd2813: data <= 8'hFF;
            13'd2814: data <= 8'h80;
            13'd2815: data <= 8'h00;
            13'd2816: data <= 8'h00;
            13'd2817: data <= 8'h00;
            13'd2818: data <= 8'h00;
            13'd2819: data <= 8'h00;
            13'd2820: data <= 8'h00;
            13'd2821: data <= 8'h00;
            13'd2822: data <= 8'h00;
            13'd2823: data <= 8'h00;
            13'd2824: data <= 8'h00;
            13'd2825: data <= 8'h03;
            13'd2826: data <= 8'hFF;
            13'd2827: data <= 8'hFF;
            13'd2828: data <= 8'hFF;
            13'd2829: data <= 8'hF8;
            13'd2830: data <= 8'h70;
            13'd2831: data <= 8'hFF;
            13'd2832: data <= 8'hE3;
            13'd2833: data <= 8'hFF;
            13'd2834: data <= 8'hFF;
            13'd2835: data <= 8'hFF;
            13'd2836: data <= 8'hFF;
            13'd2837: data <= 8'hFF;
            13'd2838: data <= 8'hFF;
            13'd2839: data <= 8'hFF;
            13'd2840: data <= 8'hFF;
            13'd2841: data <= 8'hFF;
            13'd2842: data <= 8'h01;
            13'd2843: data <= 8'hFF;
            13'd2844: data <= 8'h80;
            13'd2845: data <= 8'h00;
            13'd2846: data <= 8'h00;
            13'd2847: data <= 8'h00;
            13'd2848: data <= 8'h00;
            13'd2849: data <= 8'h00;
            13'd2850: data <= 8'h00;
            13'd2851: data <= 8'h00;
            13'd2852: data <= 8'h00;
            13'd2853: data <= 8'h00;
            13'd2854: data <= 8'h00;
            13'd2855: data <= 8'h03;
            13'd2856: data <= 8'hFF;
            13'd2857: data <= 8'hFF;
            13'd2858: data <= 8'hFF;
            13'd2859: data <= 8'hF0;
            13'd2860: data <= 8'h78;
            13'd2861: data <= 8'hFF;
            13'd2862: data <= 8'hE1;
            13'd2863: data <= 8'hFF;
            13'd2864: data <= 8'hFF;
            13'd2865: data <= 8'hFF;
            13'd2866: data <= 8'hFF;
            13'd2867: data <= 8'hFF;
            13'd2868: data <= 8'hFF;
            13'd2869: data <= 8'hFF;
            13'd2870: data <= 8'hFF;
            13'd2871: data <= 8'hFF;
            13'd2872: data <= 8'h01;
            13'd2873: data <= 8'hFF;
            13'd2874: data <= 8'h80;
            13'd2875: data <= 8'h00;
            13'd2876: data <= 8'h00;
            13'd2877: data <= 8'h00;
            13'd2878: data <= 8'h00;
            13'd2879: data <= 8'h00;
            13'd2880: data <= 8'h00;
            13'd2881: data <= 8'h00;
            13'd2882: data <= 8'h00;
            13'd2883: data <= 8'h00;
            13'd2884: data <= 8'h00;
            13'd2885: data <= 8'h03;
            13'd2886: data <= 8'hFF;
            13'd2887: data <= 8'hFF;
            13'd2888: data <= 8'hFF;
            13'd2889: data <= 8'hF0;
            13'd2890: data <= 8'h78;
            13'd2891: data <= 8'h7F;
            13'd2892: data <= 8'hE0;
            13'd2893: data <= 8'hFF;
            13'd2894: data <= 8'hFF;
            13'd2895: data <= 8'hFF;
            13'd2896: data <= 8'hFF;
            13'd2897: data <= 8'hFF;
            13'd2898: data <= 8'hFF;
            13'd2899: data <= 8'hFF;
            13'd2900: data <= 8'hFF;
            13'd2901: data <= 8'hFF;
            13'd2902: data <= 8'h80;
            13'd2903: data <= 8'hFF;
            13'd2904: data <= 8'h80;
            13'd2905: data <= 8'h00;
            13'd2906: data <= 8'h00;
            13'd2907: data <= 8'h00;
            13'd2908: data <= 8'h00;
            13'd2909: data <= 8'h00;
            13'd2910: data <= 8'h00;
            13'd2911: data <= 8'h00;
            13'd2912: data <= 8'h00;
            13'd2913: data <= 8'h00;
            13'd2914: data <= 8'h00;
            13'd2915: data <= 8'h03;
            13'd2916: data <= 8'hFF;
            13'd2917: data <= 8'hFF;
            13'd2918: data <= 8'hFF;
            13'd2919: data <= 8'hF0;
            13'd2920: data <= 8'h78;
            13'd2921: data <= 8'h7F;
            13'd2922: data <= 8'hE0;
            13'd2923: data <= 8'h7F;
            13'd2924: data <= 8'hFF;
            13'd2925: data <= 8'hFF;
            13'd2926: data <= 8'hFF;
            13'd2927: data <= 8'hFF;
            13'd2928: data <= 8'hFF;
            13'd2929: data <= 8'hFF;
            13'd2930: data <= 8'hFF;
            13'd2931: data <= 8'hFF;
            13'd2932: data <= 8'h80;
            13'd2933: data <= 8'hFF;
            13'd2934: data <= 8'h80;
            13'd2935: data <= 8'h00;
            13'd2936: data <= 8'h00;
            13'd2937: data <= 8'h00;
            13'd2938: data <= 8'h00;
            13'd2939: data <= 8'h00;
            13'd2940: data <= 8'h00;
            13'd2941: data <= 8'h00;
            13'd2942: data <= 8'h00;
            13'd2943: data <= 8'h00;
            13'd2944: data <= 8'h00;
            13'd2945: data <= 8'h03;
            13'd2946: data <= 8'hFF;
            13'd2947: data <= 8'hFF;
            13'd2948: data <= 8'hFF;
            13'd2949: data <= 8'hF0;
            13'd2950: data <= 8'h7C;
            13'd2951: data <= 8'h3F;
            13'd2952: data <= 8'hF0;
            13'd2953: data <= 8'h3F;
            13'd2954: data <= 8'hFF;
            13'd2955: data <= 8'hFF;
            13'd2956: data <= 8'hF0;
            13'd2957: data <= 8'h7F;
            13'd2958: data <= 8'hFF;
            13'd2959: data <= 8'hFF;
            13'd2960: data <= 8'hFF;
            13'd2961: data <= 8'hFF;
            13'd2962: data <= 8'hC0;
            13'd2963: data <= 8'h7F;
            13'd2964: data <= 8'h80;
            13'd2965: data <= 8'h00;
            13'd2966: data <= 8'h00;
            13'd2967: data <= 8'h00;
            13'd2968: data <= 8'h00;
            13'd2969: data <= 8'h00;
            13'd2970: data <= 8'h00;
            13'd2971: data <= 8'h00;
            13'd2972: data <= 8'h00;
            13'd2973: data <= 8'h00;
            13'd2974: data <= 8'h00;
            13'd2975: data <= 8'h03;
            13'd2976: data <= 8'hFF;
            13'd2977: data <= 8'hFF;
            13'd2978: data <= 8'hFF;
            13'd2979: data <= 8'hF8;
            13'd2980: data <= 8'h7C;
            13'd2981: data <= 8'h3F;
            13'd2982: data <= 8'hF8;
            13'd2983: data <= 8'h0F;
            13'd2984: data <= 8'hFF;
            13'd2985: data <= 8'hFF;
            13'd2986: data <= 8'hE0;
            13'd2987: data <= 8'h7F;
            13'd2988: data <= 8'hFF;
            13'd2989: data <= 8'hFF;
            13'd2990: data <= 8'hFF;
            13'd2991: data <= 8'hFF;
            13'd2992: data <= 8'hC0;
            13'd2993: data <= 8'h7F;
            13'd2994: data <= 8'h80;
            13'd2995: data <= 8'h00;
            13'd2996: data <= 8'h00;
            13'd2997: data <= 8'h00;
            13'd2998: data <= 8'h00;
            13'd2999: data <= 8'h00;
            13'd3000: data <= 8'h00;
            13'd3001: data <= 8'h00;
            13'd3002: data <= 8'h00;
            13'd3003: data <= 8'h00;
            13'd3004: data <= 8'h00;
            13'd3005: data <= 8'h03;
            13'd3006: data <= 8'hFF;
            13'd3007: data <= 8'hFF;
            13'd3008: data <= 8'hFF;
            13'd3009: data <= 8'hF8;
            13'd3010: data <= 8'h7C;
            13'd3011: data <= 8'h3F;
            13'd3012: data <= 8'hFC;
            13'd3013: data <= 8'h03;
            13'd3014: data <= 8'hFF;
            13'd3015: data <= 8'hFF;
            13'd3016: data <= 8'hC0;
            13'd3017: data <= 8'h7F;
            13'd3018: data <= 8'hFF;
            13'd3019: data <= 8'hFF;
            13'd3020: data <= 8'hFF;
            13'd3021: data <= 8'hFF;
            13'd3022: data <= 8'hC0;
            13'd3023: data <= 8'h7F;
            13'd3024: data <= 8'h80;
            13'd3025: data <= 8'h00;
            13'd3026: data <= 8'h00;
            13'd3027: data <= 8'h00;
            13'd3028: data <= 8'h00;
            13'd3029: data <= 8'h00;
            13'd3030: data <= 8'h00;
            13'd3031: data <= 8'h00;
            13'd3032: data <= 8'h00;
            13'd3033: data <= 8'h00;
            13'd3034: data <= 8'h00;
            13'd3035: data <= 8'h03;
            13'd3036: data <= 8'hFF;
            13'd3037: data <= 8'hFF;
            13'd3038: data <= 8'hFF;
            13'd3039: data <= 8'hFC;
            13'd3040: data <= 8'h7C;
            13'd3041: data <= 8'h3F;
            13'd3042: data <= 8'hFE;
            13'd3043: data <= 8'h00;
            13'd3044: data <= 8'hFF;
            13'd3045: data <= 8'hFF;
            13'd3046: data <= 8'h00;
            13'd3047: data <= 8'h7F;
            13'd3048: data <= 8'hFF;
            13'd3049: data <= 8'hFF;
            13'd3050: data <= 8'hFF;
            13'd3051: data <= 8'hFF;
            13'd3052: data <= 8'hE0;
            13'd3053: data <= 8'h3F;
            13'd3054: data <= 8'h80;
            13'd3055: data <= 8'h00;
            13'd3056: data <= 8'h00;
            13'd3057: data <= 8'h00;
            13'd3058: data <= 8'h00;
            13'd3059: data <= 8'h00;
            13'd3060: data <= 8'h00;
            13'd3061: data <= 8'h00;
            13'd3062: data <= 8'h00;
            13'd3063: data <= 8'h00;
            13'd3064: data <= 8'h00;
            13'd3065: data <= 8'h03;
            13'd3066: data <= 8'hFF;
            13'd3067: data <= 8'hFF;
            13'd3068: data <= 8'hFF;
            13'd3069: data <= 8'hFC;
            13'd3070: data <= 8'h7C;
            13'd3071: data <= 8'h1F;
            13'd3072: data <= 8'hFF;
            13'd3073: data <= 8'h80;
            13'd3074: data <= 8'h1F;
            13'd3075: data <= 8'hFE;
            13'd3076: data <= 8'h00;
            13'd3077: data <= 8'h7F;
            13'd3078: data <= 8'hFF;
            13'd3079: data <= 8'hFF;
            13'd3080: data <= 8'hFF;
            13'd3081: data <= 8'hFF;
            13'd3082: data <= 8'hE0;
            13'd3083: data <= 8'h3F;
            13'd3084: data <= 8'h80;
            13'd3085: data <= 8'h00;
            13'd3086: data <= 8'h00;
            13'd3087: data <= 8'h00;
            13'd3088: data <= 8'h00;
            13'd3089: data <= 8'h00;
            13'd3090: data <= 8'h00;
            13'd3091: data <= 8'h00;
            13'd3092: data <= 8'h00;
            13'd3093: data <= 8'h00;
            13'd3094: data <= 8'h00;
            13'd3095: data <= 8'h03;
            13'd3096: data <= 8'hFF;
            13'd3097: data <= 8'hFF;
            13'd3098: data <= 8'hFF;
            13'd3099: data <= 8'hF8;
            13'd3100: data <= 8'h7E;
            13'd3101: data <= 8'h1F;
            13'd3102: data <= 8'hFF;
            13'd3103: data <= 8'hC0;
            13'd3104: data <= 8'h03;
            13'd3105: data <= 8'h00;
            13'd3106: data <= 8'h00;
            13'd3107: data <= 8'hFF;
            13'd3108: data <= 8'hFF;
            13'd3109: data <= 8'hFF;
            13'd3110: data <= 8'hFF;
            13'd3111: data <= 8'hFF;
            13'd3112: data <= 8'hE0;
            13'd3113: data <= 8'h1F;
            13'd3114: data <= 8'h80;
            13'd3115: data <= 8'h00;
            13'd3116: data <= 8'h00;
            13'd3117: data <= 8'h00;
            13'd3118: data <= 8'h00;
            13'd3119: data <= 8'h00;
            13'd3120: data <= 8'h00;
            13'd3121: data <= 8'h00;
            13'd3122: data <= 8'h00;
            13'd3123: data <= 8'h00;
            13'd3124: data <= 8'h00;
            13'd3125: data <= 8'h03;
            13'd3126: data <= 8'hFF;
            13'd3127: data <= 8'hFF;
            13'd3128: data <= 8'hFF;
            13'd3129: data <= 8'hF8;
            13'd3130: data <= 8'h7E;
            13'd3131: data <= 8'h0F;
            13'd3132: data <= 8'hFF;
            13'd3133: data <= 8'hE0;
            13'd3134: data <= 8'h00;
            13'd3135: data <= 8'h00;
            13'd3136: data <= 8'h03;
            13'd3137: data <= 8'hFF;
            13'd3138: data <= 8'hFF;
            13'd3139: data <= 8'hFF;
            13'd3140: data <= 8'hFF;
            13'd3141: data <= 8'hFF;
            13'd3142: data <= 8'hE0;
            13'd3143: data <= 8'h1F;
            13'd3144: data <= 8'h80;
            13'd3145: data <= 8'h00;
            13'd3146: data <= 8'h00;
            13'd3147: data <= 8'h00;
            13'd3148: data <= 8'h00;
            13'd3149: data <= 8'h00;
            13'd3150: data <= 8'h00;
            13'd3151: data <= 8'h00;
            13'd3152: data <= 8'h00;
            13'd3153: data <= 8'h00;
            13'd3154: data <= 8'h00;
            13'd3155: data <= 8'h03;
            13'd3156: data <= 8'hFF;
            13'd3157: data <= 8'hFF;
            13'd3158: data <= 8'hFF;
            13'd3159: data <= 8'hF8;
            13'd3160: data <= 8'h7F;
            13'd3161: data <= 8'h0F;
            13'd3162: data <= 8'hFF;
            13'd3163: data <= 8'hF8;
            13'd3164: data <= 8'h00;
            13'd3165: data <= 8'h00;
            13'd3166: data <= 8'h07;
            13'd3167: data <= 8'hFF;
            13'd3168: data <= 8'hFF;
            13'd3169: data <= 8'hFF;
            13'd3170: data <= 8'hFF;
            13'd3171: data <= 8'hFF;
            13'd3172: data <= 8'hF0;
            13'd3173: data <= 8'h1F;
            13'd3174: data <= 8'h80;
            13'd3175: data <= 8'h00;
            13'd3176: data <= 8'h00;
            13'd3177: data <= 8'h00;
            13'd3178: data <= 8'h00;
            13'd3179: data <= 8'h00;
            13'd3180: data <= 8'h00;
            13'd3181: data <= 8'h00;
            13'd3182: data <= 8'h00;
            13'd3183: data <= 8'h00;
            13'd3184: data <= 8'h00;
            13'd3185: data <= 8'h03;
            13'd3186: data <= 8'hFF;
            13'd3187: data <= 8'hFF;
            13'd3188: data <= 8'hFF;
            13'd3189: data <= 8'hF8;
            13'd3190: data <= 8'h7F;
            13'd3191: data <= 8'h07;
            13'd3192: data <= 8'hFF;
            13'd3193: data <= 8'hFF;
            13'd3194: data <= 8'h00;
            13'd3195: data <= 8'h00;
            13'd3196: data <= 8'h1F;
            13'd3197: data <= 8'hFF;
            13'd3198: data <= 8'hFF;
            13'd3199: data <= 8'hFF;
            13'd3200: data <= 8'hFF;
            13'd3201: data <= 8'hFF;
            13'd3202: data <= 8'hF0;
            13'd3203: data <= 8'h1F;
            13'd3204: data <= 8'h80;
            13'd3205: data <= 8'h00;
            13'd3206: data <= 8'h00;
            13'd3207: data <= 8'h00;
            13'd3208: data <= 8'h00;
            13'd3209: data <= 8'h00;
            13'd3210: data <= 8'h00;
            13'd3211: data <= 8'h00;
            13'd3212: data <= 8'h00;
            13'd3213: data <= 8'h00;
            13'd3214: data <= 8'h00;
            13'd3215: data <= 8'h03;
            13'd3216: data <= 8'hFF;
            13'd3217: data <= 8'hFF;
            13'd3218: data <= 8'hFF;
            13'd3219: data <= 8'hF8;
            13'd3220: data <= 8'h7F;
            13'd3221: data <= 8'h87;
            13'd3222: data <= 8'hFF;
            13'd3223: data <= 8'hFF;
            13'd3224: data <= 8'hF0;
            13'd3225: data <= 8'h00;
            13'd3226: data <= 8'h7F;
            13'd3227: data <= 8'hFF;
            13'd3228: data <= 8'hFF;
            13'd3229: data <= 8'hFF;
            13'd3230: data <= 8'hFF;
            13'd3231: data <= 8'hFF;
            13'd3232: data <= 8'hF8;
            13'd3233: data <= 8'h0F;
            13'd3234: data <= 8'h80;
            13'd3235: data <= 8'h00;
            13'd3236: data <= 8'h00;
            13'd3237: data <= 8'h00;
            13'd3238: data <= 8'h00;
            13'd3239: data <= 8'h00;
            13'd3240: data <= 8'h00;
            13'd3241: data <= 8'h00;
            13'd3242: data <= 8'h00;
            13'd3243: data <= 8'h00;
            13'd3244: data <= 8'h00;
            13'd3245: data <= 8'h03;
            13'd3246: data <= 8'hFF;
            13'd3247: data <= 8'hFF;
            13'd3248: data <= 8'hFF;
            13'd3249: data <= 8'hF8;
            13'd3250: data <= 8'h7F;
            13'd3251: data <= 8'h83;
            13'd3252: data <= 8'hFF;
            13'd3253: data <= 8'hFF;
            13'd3254: data <= 8'hFE;
            13'd3255: data <= 8'h01;
            13'd3256: data <= 8'hFF;
            13'd3257: data <= 8'hFF;
            13'd3258: data <= 8'hFF;
            13'd3259: data <= 8'hFF;
            13'd3260: data <= 8'hFF;
            13'd3261: data <= 8'hFF;
            13'd3262: data <= 8'hF8;
            13'd3263: data <= 8'h0F;
            13'd3264: data <= 8'h80;
            13'd3265: data <= 8'h00;
            13'd3266: data <= 8'h00;
            13'd3267: data <= 8'h00;
            13'd3268: data <= 8'h00;
            13'd3269: data <= 8'h00;
            13'd3270: data <= 8'h00;
            13'd3271: data <= 8'h00;
            13'd3272: data <= 8'h00;
            13'd3273: data <= 8'h00;
            13'd3274: data <= 8'h00;
            13'd3275: data <= 8'h03;
            13'd3276: data <= 8'hFF;
            13'd3277: data <= 8'hFF;
            13'd3278: data <= 8'hFF;
            13'd3279: data <= 8'hF8;
            13'd3280: data <= 8'h7F;
            13'd3281: data <= 8'hC1;
            13'd3282: data <= 8'hFF;
            13'd3283: data <= 8'hFF;
            13'd3284: data <= 8'hFF;
            13'd3285: data <= 8'hFF;
            13'd3286: data <= 8'hFF;
            13'd3287: data <= 8'hFF;
            13'd3288: data <= 8'hFF;
            13'd3289: data <= 8'hFF;
            13'd3290: data <= 8'hFF;
            13'd3291: data <= 8'hFF;
            13'd3292: data <= 8'hF8;
            13'd3293: data <= 8'h0F;
            13'd3294: data <= 8'h80;
            13'd3295: data <= 8'h00;
            13'd3296: data <= 8'h00;
            13'd3297: data <= 8'h00;
            13'd3298: data <= 8'h00;
            13'd3299: data <= 8'h00;
            13'd3300: data <= 8'h00;
            13'd3301: data <= 8'h00;
            13'd3302: data <= 8'h00;
            13'd3303: data <= 8'h00;
            13'd3304: data <= 8'h00;
            13'd3305: data <= 8'h03;
            13'd3306: data <= 8'hFF;
            13'd3307: data <= 8'hFF;
            13'd3308: data <= 8'hFF;
            13'd3309: data <= 8'hF8;
            13'd3310: data <= 8'h7F;
            13'd3311: data <= 8'hC1;
            13'd3312: data <= 8'hFF;
            13'd3313: data <= 8'hFF;
            13'd3314: data <= 8'hFF;
            13'd3315: data <= 8'hFF;
            13'd3316: data <= 8'hFF;
            13'd3317: data <= 8'hFF;
            13'd3318: data <= 8'hFF;
            13'd3319: data <= 8'hFF;
            13'd3320: data <= 8'hFF;
            13'd3321: data <= 8'hFF;
            13'd3322: data <= 8'hF8;
            13'd3323: data <= 8'h07;
            13'd3324: data <= 8'h80;
            13'd3325: data <= 8'h00;
            13'd3326: data <= 8'h00;
            13'd3327: data <= 8'h00;
            13'd3328: data <= 8'h00;
            13'd3329: data <= 8'h00;
            13'd3330: data <= 8'h00;
            13'd3331: data <= 8'h00;
            13'd3332: data <= 8'h00;
            13'd3333: data <= 8'h00;
            13'd3334: data <= 8'h00;
            13'd3335: data <= 8'h03;
            13'd3336: data <= 8'hFF;
            13'd3337: data <= 8'hFF;
            13'd3338: data <= 8'hFF;
            13'd3339: data <= 8'hF8;
            13'd3340: data <= 8'h7F;
            13'd3341: data <= 8'hE0;
            13'd3342: data <= 8'hFF;
            13'd3343: data <= 8'hFF;
            13'd3344: data <= 8'hFF;
            13'd3345: data <= 8'hFF;
            13'd3346: data <= 8'hFF;
            13'd3347: data <= 8'hFF;
            13'd3348: data <= 8'hFF;
            13'd3349: data <= 8'hFF;
            13'd3350: data <= 8'hFF;
            13'd3351: data <= 8'hFF;
            13'd3352: data <= 8'hFC;
            13'd3353: data <= 8'h07;
            13'd3354: data <= 8'h80;
            13'd3355: data <= 8'h00;
            13'd3356: data <= 8'h00;
            13'd3357: data <= 8'h00;
            13'd3358: data <= 8'h00;
            13'd3359: data <= 8'h00;
            13'd3360: data <= 8'h00;
            13'd3361: data <= 8'h00;
            13'd3362: data <= 8'h00;
            13'd3363: data <= 8'h00;
            13'd3364: data <= 8'h00;
            13'd3365: data <= 8'h03;
            13'd3366: data <= 8'hFF;
            13'd3367: data <= 8'hFF;
            13'd3368: data <= 8'hFF;
            13'd3369: data <= 8'hFC;
            13'd3370: data <= 8'h7F;
            13'd3371: data <= 8'hE0;
            13'd3372: data <= 8'h7F;
            13'd3373: data <= 8'hFF;
            13'd3374: data <= 8'hFF;
            13'd3375: data <= 8'hFF;
            13'd3376: data <= 8'hFF;
            13'd3377: data <= 8'hFF;
            13'd3378: data <= 8'hFF;
            13'd3379: data <= 8'hFF;
            13'd3380: data <= 8'hFF;
            13'd3381: data <= 8'hFF;
            13'd3382: data <= 8'hFC;
            13'd3383: data <= 8'h07;
            13'd3384: data <= 8'h80;
            13'd3385: data <= 8'h00;
            13'd3386: data <= 8'h00;
            13'd3387: data <= 8'h00;
            13'd3388: data <= 8'h00;
            13'd3389: data <= 8'h00;
            13'd3390: data <= 8'h00;
            13'd3391: data <= 8'h00;
            13'd3392: data <= 8'h00;
            13'd3393: data <= 8'h00;
            13'd3394: data <= 8'h00;
            13'd3395: data <= 8'h03;
            13'd3396: data <= 8'hFF;
            13'd3397: data <= 8'hFF;
            13'd3398: data <= 8'hFF;
            13'd3399: data <= 8'hFC;
            13'd3400: data <= 8'h7F;
            13'd3401: data <= 8'hF0;
            13'd3402: data <= 8'h7F;
            13'd3403: data <= 8'hFF;
            13'd3404: data <= 8'hFF;
            13'd3405: data <= 8'hFF;
            13'd3406: data <= 8'hFF;
            13'd3407: data <= 8'hFF;
            13'd3408: data <= 8'hFF;
            13'd3409: data <= 8'hFF;
            13'd3410: data <= 8'hFF;
            13'd3411: data <= 8'hFF;
            13'd3412: data <= 8'hFC;
            13'd3413: data <= 8'h03;
            13'd3414: data <= 8'h80;
            13'd3415: data <= 8'h00;
            13'd3416: data <= 8'h00;
            13'd3417: data <= 8'h00;
            13'd3418: data <= 8'h00;
            13'd3419: data <= 8'h00;
            13'd3420: data <= 8'h00;
            13'd3421: data <= 8'h00;
            13'd3422: data <= 8'h00;
            13'd3423: data <= 8'h00;
            13'd3424: data <= 8'h00;
            13'd3425: data <= 8'h03;
            13'd3426: data <= 8'hFF;
            13'd3427: data <= 8'hFF;
            13'd3428: data <= 8'hFF;
            13'd3429: data <= 8'hFC;
            13'd3430: data <= 8'h7F;
            13'd3431: data <= 8'hF8;
            13'd3432: data <= 8'h3F;
            13'd3433: data <= 8'hFF;
            13'd3434: data <= 8'hFF;
            13'd3435: data <= 8'hFF;
            13'd3436: data <= 8'hFF;
            13'd3437: data <= 8'hFF;
            13'd3438: data <= 8'hFF;
            13'd3439: data <= 8'hFF;
            13'd3440: data <= 8'hFF;
            13'd3441: data <= 8'hFF;
            13'd3442: data <= 8'hFE;
            13'd3443: data <= 8'h03;
            13'd3444: data <= 8'h80;
            13'd3445: data <= 8'h00;
            13'd3446: data <= 8'h00;
            13'd3447: data <= 8'h00;
            13'd3448: data <= 8'h00;
            13'd3449: data <= 8'h00;
            13'd3450: data <= 8'h00;
            13'd3451: data <= 8'h00;
            13'd3452: data <= 8'h00;
            13'd3453: data <= 8'h00;
            13'd3454: data <= 8'h00;
            13'd3455: data <= 8'h03;
            13'd3456: data <= 8'hFF;
            13'd3457: data <= 8'hFF;
            13'd3458: data <= 8'hFF;
            13'd3459: data <= 8'hFC;
            13'd3460: data <= 8'h7F;
            13'd3461: data <= 8'hFC;
            13'd3462: data <= 8'h1F;
            13'd3463: data <= 8'hFF;
            13'd3464: data <= 8'hFF;
            13'd3465: data <= 8'hFF;
            13'd3466: data <= 8'hFF;
            13'd3467: data <= 8'hFF;
            13'd3468: data <= 8'hFF;
            13'd3469: data <= 8'hFF;
            13'd3470: data <= 8'hFF;
            13'd3471: data <= 8'hFF;
            13'd3472: data <= 8'hFE;
            13'd3473: data <= 8'h03;
            13'd3474: data <= 8'h80;
            13'd3475: data <= 8'h00;
            13'd3476: data <= 8'h00;
            13'd3477: data <= 8'h00;
            13'd3478: data <= 8'h00;
            13'd3479: data <= 8'h00;
            13'd3480: data <= 8'h00;
            13'd3481: data <= 8'h00;
            13'd3482: data <= 8'h00;
            13'd3483: data <= 8'h00;
            13'd3484: data <= 8'h00;
            13'd3485: data <= 8'h03;
            13'd3486: data <= 8'hFF;
            13'd3487: data <= 8'hFF;
            13'd3488: data <= 8'hFF;
            13'd3489: data <= 8'hFC;
            13'd3490: data <= 8'h7F;
            13'd3491: data <= 8'hFC;
            13'd3492: data <= 8'h0F;
            13'd3493: data <= 8'hFF;
            13'd3494: data <= 8'hFF;
            13'd3495: data <= 8'hFF;
            13'd3496: data <= 8'hFF;
            13'd3497: data <= 8'hFF;
            13'd3498: data <= 8'hFF;
            13'd3499: data <= 8'hFF;
            13'd3500: data <= 8'hFF;
            13'd3501: data <= 8'hFF;
            13'd3502: data <= 8'hFE;
            13'd3503: data <= 8'h03;
            13'd3504: data <= 8'h80;
            13'd3505: data <= 8'h00;
            13'd3506: data <= 8'h00;
            13'd3507: data <= 8'h00;
            13'd3508: data <= 8'h00;
            13'd3509: data <= 8'h00;
            13'd3510: data <= 8'h00;
            13'd3511: data <= 8'h00;
            13'd3512: data <= 8'h00;
            13'd3513: data <= 8'h00;
            13'd3514: data <= 8'h00;
            13'd3515: data <= 8'h03;
            13'd3516: data <= 8'hFF;
            13'd3517: data <= 8'hFF;
            13'd3518: data <= 8'hFF;
            13'd3519: data <= 8'hFC;
            13'd3520: data <= 8'h7F;
            13'd3521: data <= 8'hFE;
            13'd3522: data <= 8'h07;
            13'd3523: data <= 8'hFF;
            13'd3524: data <= 8'hFF;
            13'd3525: data <= 8'hFF;
            13'd3526: data <= 8'hFF;
            13'd3527: data <= 8'hFF;
            13'd3528: data <= 8'hFF;
            13'd3529: data <= 8'hFF;
            13'd3530: data <= 8'hFF;
            13'd3531: data <= 8'hFF;
            13'd3532: data <= 8'hFF;
            13'd3533: data <= 8'h03;
            13'd3534: data <= 8'h80;
            13'd3535: data <= 8'h00;
            13'd3536: data <= 8'h00;
            13'd3537: data <= 8'h00;
            13'd3538: data <= 8'h00;
            13'd3539: data <= 8'h00;
            13'd3540: data <= 8'h00;
            13'd3541: data <= 8'h00;
            13'd3542: data <= 8'h00;
            13'd3543: data <= 8'h00;
            13'd3544: data <= 8'h00;
            13'd3545: data <= 8'h03;
            13'd3546: data <= 8'hFF;
            13'd3547: data <= 8'hFF;
            13'd3548: data <= 8'hFF;
            13'd3549: data <= 8'hFC;
            13'd3550: data <= 8'h7F;
            13'd3551: data <= 8'hFF;
            13'd3552: data <= 8'h03;
            13'd3553: data <= 8'hFF;
            13'd3554: data <= 8'hFF;
            13'd3555: data <= 8'hFF;
            13'd3556: data <= 8'hFF;
            13'd3557: data <= 8'hFF;
            13'd3558: data <= 8'hFF;
            13'd3559: data <= 8'hFF;
            13'd3560: data <= 8'hFF;
            13'd3561: data <= 8'hFF;
            13'd3562: data <= 8'hFF;
            13'd3563: data <= 8'h01;
            13'd3564: data <= 8'h80;
            13'd3565: data <= 8'h00;
            13'd3566: data <= 8'h00;
            13'd3567: data <= 8'h00;
            13'd3568: data <= 8'h00;
            13'd3569: data <= 8'h00;
            13'd3570: data <= 8'h00;
            13'd3571: data <= 8'h00;
            13'd3572: data <= 8'h00;
            13'd3573: data <= 8'h00;
            13'd3574: data <= 8'h00;
            13'd3575: data <= 8'h03;
            13'd3576: data <= 8'hFF;
            13'd3577: data <= 8'hFF;
            13'd3578: data <= 8'hFF;
            13'd3579: data <= 8'hFC;
            13'd3580: data <= 8'h7F;
            13'd3581: data <= 8'hFF;
            13'd3582: data <= 8'h81;
            13'd3583: data <= 8'hFF;
            13'd3584: data <= 8'hFF;
            13'd3585: data <= 8'hFF;
            13'd3586: data <= 8'hFF;
            13'd3587: data <= 8'hFF;
            13'd3588: data <= 8'hFF;
            13'd3589: data <= 8'hFF;
            13'd3590: data <= 8'hFF;
            13'd3591: data <= 8'hFF;
            13'd3592: data <= 8'hFF;
            13'd3593: data <= 8'h81;
            13'd3594: data <= 8'h80;
            13'd3595: data <= 8'h00;
            13'd3596: data <= 8'h00;
            13'd3597: data <= 8'h00;
            13'd3598: data <= 8'h00;
            13'd3599: data <= 8'h00;
            13'd3600: data <= 8'h00;
            13'd3601: data <= 8'h00;
            13'd3602: data <= 8'h00;
            13'd3603: data <= 8'h00;
            13'd3604: data <= 8'h00;
            13'd3605: data <= 8'h03;
            13'd3606: data <= 8'hFF;
            13'd3607: data <= 8'hFF;
            13'd3608: data <= 8'hFF;
            13'd3609: data <= 8'hFC;
            13'd3610: data <= 8'h7F;
            13'd3611: data <= 8'hFF;
            13'd3612: data <= 8'hC1;
            13'd3613: data <= 8'hFF;
            13'd3614: data <= 8'hFF;
            13'd3615: data <= 8'hFF;
            13'd3616: data <= 8'hFF;
            13'd3617: data <= 8'hFF;
            13'd3618: data <= 8'hFF;
            13'd3619: data <= 8'hFF;
            13'd3620: data <= 8'hFF;
            13'd3621: data <= 8'hFF;
            13'd3622: data <= 8'hFF;
            13'd3623: data <= 8'h81;
            13'd3624: data <= 8'h80;
            13'd3625: data <= 8'h00;
            13'd3626: data <= 8'h00;
            13'd3627: data <= 8'h00;
            13'd3628: data <= 8'h00;
            13'd3629: data <= 8'h00;
            13'd3630: data <= 8'h00;
            13'd3631: data <= 8'h00;
            13'd3632: data <= 8'h00;
            13'd3633: data <= 8'h00;
            13'd3634: data <= 8'h00;
            13'd3635: data <= 8'h03;
            13'd3636: data <= 8'hFF;
            13'd3637: data <= 8'hFF;
            13'd3638: data <= 8'hFF;
            13'd3639: data <= 8'hF8;
            13'd3640: data <= 8'h7F;
            13'd3641: data <= 8'hFF;
            13'd3642: data <= 8'hE0;
            13'd3643: data <= 8'h7F;
            13'd3644: data <= 8'hFF;
            13'd3645: data <= 8'hFF;
            13'd3646: data <= 8'hFF;
            13'd3647: data <= 8'hFF;
            13'd3648: data <= 8'hFF;
            13'd3649: data <= 8'hFF;
            13'd3650: data <= 8'hFF;
            13'd3651: data <= 8'hFF;
            13'd3652: data <= 8'hFF;
            13'd3653: data <= 8'h81;
            13'd3654: data <= 8'h80;
            13'd3655: data <= 8'h00;
            13'd3656: data <= 8'h00;
            13'd3657: data <= 8'h00;
            13'd3658: data <= 8'h00;
            13'd3659: data <= 8'h00;
            13'd3660: data <= 8'h00;
            13'd3661: data <= 8'h00;
            13'd3662: data <= 8'h00;
            13'd3663: data <= 8'h00;
            13'd3664: data <= 8'h00;
            13'd3665: data <= 8'h03;
            13'd3666: data <= 8'hFF;
            13'd3667: data <= 8'hFF;
            13'd3668: data <= 8'hFF;
            13'd3669: data <= 8'hF0;
            13'd3670: data <= 8'h7F;
            13'd3671: data <= 8'hFF;
            13'd3672: data <= 8'hF0;
            13'd3673: data <= 8'h3F;
            13'd3674: data <= 8'hFF;
            13'd3675: data <= 8'hFF;
            13'd3676: data <= 8'hFF;
            13'd3677: data <= 8'hFF;
            13'd3678: data <= 8'hFF;
            13'd3679: data <= 8'hFF;
            13'd3680: data <= 8'hFF;
            13'd3681: data <= 8'hFF;
            13'd3682: data <= 8'hFF;
            13'd3683: data <= 8'h80;
            13'd3684: data <= 8'h80;
            13'd3685: data <= 8'h00;
            13'd3686: data <= 8'h00;
            13'd3687: data <= 8'h00;
            13'd3688: data <= 8'h00;
            13'd3689: data <= 8'h00;
            13'd3690: data <= 8'h00;
            13'd3691: data <= 8'h00;
            13'd3692: data <= 8'h00;
            13'd3693: data <= 8'h00;
            13'd3694: data <= 8'h00;
            13'd3695: data <= 8'h03;
            13'd3696: data <= 8'hFF;
            13'd3697: data <= 8'hFF;
            13'd3698: data <= 8'hFF;
            13'd3699: data <= 8'hF0;
            13'd3700: data <= 8'h7F;
            13'd3701: data <= 8'hFF;
            13'd3702: data <= 8'hF0;
            13'd3703: data <= 8'h1F;
            13'd3704: data <= 8'hFF;
            13'd3705: data <= 8'hFF;
            13'd3706: data <= 8'hFF;
            13'd3707: data <= 8'hFF;
            13'd3708: data <= 8'hFF;
            13'd3709: data <= 8'hFF;
            13'd3710: data <= 8'hFF;
            13'd3711: data <= 8'hFF;
            13'd3712: data <= 8'hFF;
            13'd3713: data <= 8'h80;
            13'd3714: data <= 8'h80;
            13'd3715: data <= 8'h00;
            13'd3716: data <= 8'h00;
            13'd3717: data <= 8'h00;
            13'd3718: data <= 8'h00;
            13'd3719: data <= 8'h00;
            13'd3720: data <= 8'h00;
            13'd3721: data <= 8'h00;
            13'd3722: data <= 8'h00;
            13'd3723: data <= 8'h00;
            13'd3724: data <= 8'h00;
            13'd3725: data <= 8'h03;
            13'd3726: data <= 8'hFF;
            13'd3727: data <= 8'hFF;
            13'd3728: data <= 8'hFF;
            13'd3729: data <= 8'hF0;
            13'd3730: data <= 8'h3F;
            13'd3731: data <= 8'hFF;
            13'd3732: data <= 8'hF8;
            13'd3733: data <= 8'h07;
            13'd3734: data <= 8'hFF;
            13'd3735: data <= 8'hFF;
            13'd3736: data <= 8'hFF;
            13'd3737: data <= 8'hFF;
            13'd3738: data <= 8'hFF;
            13'd3739: data <= 8'hFF;
            13'd3740: data <= 8'hFF;
            13'd3741: data <= 8'hFF;
            13'd3742: data <= 8'hFF;
            13'd3743: data <= 8'h80;
            13'd3744: data <= 8'h80;
            13'd3745: data <= 8'h00;
            13'd3746: data <= 8'h00;
            13'd3747: data <= 8'h00;
            13'd3748: data <= 8'h00;
            13'd3749: data <= 8'h00;
            13'd3750: data <= 8'h00;
            13'd3751: data <= 8'h00;
            13'd3752: data <= 8'h00;
            13'd3753: data <= 8'h00;
            13'd3754: data <= 8'h00;
            13'd3755: data <= 8'h03;
            13'd3756: data <= 8'hFF;
            13'd3757: data <= 8'hFF;
            13'd3758: data <= 8'hFF;
            13'd3759: data <= 8'hF8;
            13'd3760: data <= 8'h3F;
            13'd3761: data <= 8'hFF;
            13'd3762: data <= 8'hFE;
            13'd3763: data <= 8'h01;
            13'd3764: data <= 8'hFF;
            13'd3765: data <= 8'hFF;
            13'd3766: data <= 8'hFF;
            13'd3767: data <= 8'hFF;
            13'd3768: data <= 8'hFF;
            13'd3769: data <= 8'hFF;
            13'd3770: data <= 8'hFF;
            13'd3771: data <= 8'hFF;
            13'd3772: data <= 8'hFF;
            13'd3773: data <= 8'hC0;
            13'd3774: data <= 8'h00;
            13'd3775: data <= 8'h00;
            13'd3776: data <= 8'h00;
            13'd3777: data <= 8'h00;
            13'd3778: data <= 8'h00;
            13'd3779: data <= 8'h00;
            13'd3780: data <= 8'h00;
            13'd3781: data <= 8'h00;
            13'd3782: data <= 8'h00;
            13'd3783: data <= 8'h00;
            13'd3784: data <= 8'h00;
            13'd3785: data <= 8'h03;
            13'd3786: data <= 8'hFF;
            13'd3787: data <= 8'hFF;
            13'd3788: data <= 8'hFF;
            13'd3789: data <= 8'hF8;
            13'd3790: data <= 8'h3F;
            13'd3791: data <= 8'hFF;
            13'd3792: data <= 8'hFF;
            13'd3793: data <= 8'h00;
            13'd3794: data <= 8'hFF;
            13'd3795: data <= 8'hFF;
            13'd3796: data <= 8'hFF;
            13'd3797: data <= 8'hFF;
            13'd3798: data <= 8'hFF;
            13'd3799: data <= 8'hFF;
            13'd3800: data <= 8'hFF;
            13'd3801: data <= 8'hFF;
            13'd3802: data <= 8'hFF;
            13'd3803: data <= 8'hC0;
            13'd3804: data <= 8'h00;
            13'd3805: data <= 8'h00;
            13'd3806: data <= 8'h00;
            13'd3807: data <= 8'h00;
            13'd3808: data <= 8'h00;
            13'd3809: data <= 8'h00;
            13'd3810: data <= 8'h00;
            13'd3811: data <= 8'h00;
            13'd3812: data <= 8'h00;
            13'd3813: data <= 8'h00;
            13'd3814: data <= 8'h00;
            13'd3815: data <= 8'h03;
            13'd3816: data <= 8'hFF;
            13'd3817: data <= 8'hFF;
            13'd3818: data <= 8'hFF;
            13'd3819: data <= 8'hF8;
            13'd3820: data <= 8'h7F;
            13'd3821: data <= 8'hFF;
            13'd3822: data <= 8'hFF;
            13'd3823: data <= 8'h80;
            13'd3824: data <= 8'h1F;
            13'd3825: data <= 8'hFF;
            13'd3826: data <= 8'hFF;
            13'd3827: data <= 8'hFF;
            13'd3828: data <= 8'hFF;
            13'd3829: data <= 8'hFF;
            13'd3830: data <= 8'hFF;
            13'd3831: data <= 8'hFF;
            13'd3832: data <= 8'hFF;
            13'd3833: data <= 8'hC0;
            13'd3834: data <= 8'h00;
            13'd3835: data <= 8'h00;
            13'd3836: data <= 8'h00;
            13'd3837: data <= 8'h00;
            13'd3838: data <= 8'h00;
            13'd3839: data <= 8'h00;
            13'd3840: data <= 8'h00;
            13'd3841: data <= 8'h00;
            13'd3842: data <= 8'h00;
            13'd3843: data <= 8'h00;
            13'd3844: data <= 8'h00;
            13'd3845: data <= 8'h03;
            13'd3846: data <= 8'hFF;
            13'd3847: data <= 8'hFF;
            13'd3848: data <= 8'hFF;
            13'd3849: data <= 8'hF8;
            13'd3850: data <= 8'h7F;
            13'd3851: data <= 8'hFF;
            13'd3852: data <= 8'hFF;
            13'd3853: data <= 8'hC0;
            13'd3854: data <= 8'h07;
            13'd3855: data <= 8'hFF;
            13'd3856: data <= 8'hFF;
            13'd3857: data <= 8'hFF;
            13'd3858: data <= 8'hFF;
            13'd3859: data <= 8'hFF;
            13'd3860: data <= 8'hFF;
            13'd3861: data <= 8'hFF;
            13'd3862: data <= 8'hFF;
            13'd3863: data <= 8'hC0;
            13'd3864: data <= 8'h00;
            13'd3865: data <= 8'h00;
            13'd3866: data <= 8'h00;
            13'd3867: data <= 8'h00;
            13'd3868: data <= 8'h00;
            13'd3869: data <= 8'h00;
            13'd3870: data <= 8'h00;
            13'd3871: data <= 8'h00;
            13'd3872: data <= 8'h00;
            13'd3873: data <= 8'h00;
            13'd3874: data <= 8'h00;
            13'd3875: data <= 8'h03;
            13'd3876: data <= 8'hFF;
            13'd3877: data <= 8'hFF;
            13'd3878: data <= 8'hFF;
            13'd3879: data <= 8'hF8;
            13'd3880: data <= 8'h7F;
            13'd3881: data <= 8'hFF;
            13'd3882: data <= 8'hFF;
            13'd3883: data <= 8'hE0;
            13'd3884: data <= 8'h01;
            13'd3885: data <= 8'hFF;
            13'd3886: data <= 8'hFF;
            13'd3887: data <= 8'hFF;
            13'd3888: data <= 8'hFF;
            13'd3889: data <= 8'hFF;
            13'd3890: data <= 8'hFF;
            13'd3891: data <= 8'hFF;
            13'd3892: data <= 8'hFF;
            13'd3893: data <= 8'hC0;
            13'd3894: data <= 8'h00;
            13'd3895: data <= 8'h00;
            13'd3896: data <= 8'h00;
            13'd3897: data <= 8'h00;
            13'd3898: data <= 8'h00;
            13'd3899: data <= 8'h00;
            13'd3900: data <= 8'h00;
            13'd3901: data <= 8'h00;
            13'd3902: data <= 8'h00;
            13'd3903: data <= 8'h00;
            13'd3904: data <= 8'h00;
            13'd3905: data <= 8'h03;
            13'd3906: data <= 8'hFF;
            13'd3907: data <= 8'hFF;
            13'd3908: data <= 8'hFF;
            13'd3909: data <= 8'hF8;
            13'd3910: data <= 8'h7F;
            13'd3911: data <= 8'hFF;
            13'd3912: data <= 8'hFF;
            13'd3913: data <= 8'hF8;
            13'd3914: data <= 8'h00;
            13'd3915: data <= 8'h7F;
            13'd3916: data <= 8'hFC;
            13'd3917: data <= 8'h7F;
            13'd3918: data <= 8'hFF;
            13'd3919: data <= 8'hFF;
            13'd3920: data <= 8'hFF;
            13'd3921: data <= 8'hFF;
            13'd3922: data <= 8'hFF;
            13'd3923: data <= 8'hE0;
            13'd3924: data <= 8'h00;
            13'd3925: data <= 8'h00;
            13'd3926: data <= 8'h00;
            13'd3927: data <= 8'h00;
            13'd3928: data <= 8'h00;
            13'd3929: data <= 8'h00;
            13'd3930: data <= 8'h00;
            13'd3931: data <= 8'h00;
            13'd3932: data <= 8'h00;
            13'd3933: data <= 8'h00;
            13'd3934: data <= 8'h00;
            13'd3935: data <= 8'h03;
            13'd3936: data <= 8'hFF;
            13'd3937: data <= 8'hFF;
            13'd3938: data <= 8'hFF;
            13'd3939: data <= 8'hF8;
            13'd3940: data <= 8'h7F;
            13'd3941: data <= 8'hFF;
            13'd3942: data <= 8'hFF;
            13'd3943: data <= 8'hFC;
            13'd3944: data <= 8'h00;
            13'd3945: data <= 8'h00;
            13'd3946: data <= 8'hC0;
            13'd3947: data <= 8'h3F;
            13'd3948: data <= 8'hFF;
            13'd3949: data <= 8'hFF;
            13'd3950: data <= 8'hFF;
            13'd3951: data <= 8'hFF;
            13'd3952: data <= 8'hFF;
            13'd3953: data <= 8'hE0;
            13'd3954: data <= 8'h00;
            13'd3955: data <= 8'h00;
            13'd3956: data <= 8'h00;
            13'd3957: data <= 8'h00;
            13'd3958: data <= 8'h00;
            13'd3959: data <= 8'h00;
            13'd3960: data <= 8'h00;
            13'd3961: data <= 8'h00;
            13'd3962: data <= 8'h00;
            13'd3963: data <= 8'h00;
            13'd3964: data <= 8'h00;
            13'd3965: data <= 8'h03;
            13'd3966: data <= 8'hFF;
            13'd3967: data <= 8'hFF;
            13'd3968: data <= 8'hFF;
            13'd3969: data <= 8'hF0;
            13'd3970: data <= 8'h7F;
            13'd3971: data <= 8'hFF;
            13'd3972: data <= 8'hFF;
            13'd3973: data <= 8'hFF;
            13'd3974: data <= 8'h00;
            13'd3975: data <= 8'h00;
            13'd3976: data <= 8'h00;
            13'd3977: data <= 8'h1F;
            13'd3978: data <= 8'hFF;
            13'd3979: data <= 8'hFF;
            13'd3980: data <= 8'hFF;
            13'd3981: data <= 8'hFF;
            13'd3982: data <= 8'hFF;
            13'd3983: data <= 8'hE0;
            13'd3984: data <= 8'h00;
            13'd3985: data <= 8'h00;
            13'd3986: data <= 8'h00;
            13'd3987: data <= 8'h00;
            13'd3988: data <= 8'h00;
            13'd3989: data <= 8'h00;
            13'd3990: data <= 8'h00;
            13'd3991: data <= 8'h00;
            13'd3992: data <= 8'h00;
            13'd3993: data <= 8'h00;
            13'd3994: data <= 8'h00;
            13'd3995: data <= 8'h03;
            13'd3996: data <= 8'hFF;
            13'd3997: data <= 8'hFF;
            13'd3998: data <= 8'hFF;
            13'd3999: data <= 8'hF0;
            13'd4000: data <= 8'h7F;
            13'd4001: data <= 8'hFF;
            13'd4002: data <= 8'hFF;
            13'd4003: data <= 8'hFF;
            13'd4004: data <= 8'hC0;
            13'd4005: data <= 8'h00;
            13'd4006: data <= 8'h00;
            13'd4007: data <= 8'h3F;
            13'd4008: data <= 8'hFF;
            13'd4009: data <= 8'hFF;
            13'd4010: data <= 8'hFF;
            13'd4011: data <= 8'hFF;
            13'd4012: data <= 8'hFF;
            13'd4013: data <= 8'hE0;
            13'd4014: data <= 8'h00;
            13'd4015: data <= 8'h00;
            13'd4016: data <= 8'h00;
            13'd4017: data <= 8'h00;
            13'd4018: data <= 8'h00;
            13'd4019: data <= 8'h00;
            13'd4020: data <= 8'h00;
            13'd4021: data <= 8'h00;
            13'd4022: data <= 8'h00;
            13'd4023: data <= 8'h00;
            13'd4024: data <= 8'h00;
            13'd4025: data <= 8'h03;
            13'd4026: data <= 8'hFF;
            13'd4027: data <= 8'hFF;
            13'd4028: data <= 8'hFF;
            13'd4029: data <= 8'hF0;
            13'd4030: data <= 8'h7F;
            13'd4031: data <= 8'hFF;
            13'd4032: data <= 8'hFF;
            13'd4033: data <= 8'hFF;
            13'd4034: data <= 8'hF0;
            13'd4035: data <= 8'h00;
            13'd4036: data <= 8'h00;
            13'd4037: data <= 8'h3F;
            13'd4038: data <= 8'hFF;
            13'd4039: data <= 8'hFF;
            13'd4040: data <= 8'hFF;
            13'd4041: data <= 8'hFF;
            13'd4042: data <= 8'hFF;
            13'd4043: data <= 8'hE0;
            13'd4044: data <= 8'h00;
            13'd4045: data <= 8'h00;
            13'd4046: data <= 8'h00;
            13'd4047: data <= 8'h00;
            13'd4048: data <= 8'h00;
            13'd4049: data <= 8'h00;
            13'd4050: data <= 8'h00;
            13'd4051: data <= 8'h00;
            13'd4052: data <= 8'h00;
            13'd4053: data <= 8'h00;
            13'd4054: data <= 8'h00;
            13'd4055: data <= 8'h03;
            13'd4056: data <= 8'hFF;
            13'd4057: data <= 8'hFF;
            13'd4058: data <= 8'hFF;
            13'd4059: data <= 8'hF0;
            13'd4060: data <= 8'h7F;
            13'd4061: data <= 8'hFF;
            13'd4062: data <= 8'hFF;
            13'd4063: data <= 8'hFF;
            13'd4064: data <= 8'hF8;
            13'd4065: data <= 8'h00;
            13'd4066: data <= 8'h00;
            13'd4067: data <= 8'h7F;
            13'd4068: data <= 8'hFF;
            13'd4069: data <= 8'hFF;
            13'd4070: data <= 8'hFF;
            13'd4071: data <= 8'hFF;
            13'd4072: data <= 8'hFF;
            13'd4073: data <= 8'hE0;
            13'd4074: data <= 8'h00;
            13'd4075: data <= 8'h00;
            13'd4076: data <= 8'h00;
            13'd4077: data <= 8'h00;
            13'd4078: data <= 8'h00;
            13'd4079: data <= 8'h00;
            13'd4080: data <= 8'h00;
            13'd4081: data <= 8'h00;
            13'd4082: data <= 8'h00;
            13'd4083: data <= 8'h00;
            13'd4084: data <= 8'h00;
            13'd4085: data <= 8'h03;
            13'd4086: data <= 8'hFF;
            13'd4087: data <= 8'hFF;
            13'd4088: data <= 8'hFF;
            13'd4089: data <= 8'hF0;
            13'd4090: data <= 8'h7F;
            13'd4091: data <= 8'hFF;
            13'd4092: data <= 8'hFF;
            13'd4093: data <= 8'hFF;
            13'd4094: data <= 8'hFF;
            13'd4095: data <= 8'hC0;
            13'd4096: data <= 8'h03;
            13'd4097: data <= 8'hFF;
            13'd4098: data <= 8'hFF;
            13'd4099: data <= 8'hFF;
            13'd4100: data <= 8'hFF;
            13'd4101: data <= 8'hFF;
            13'd4102: data <= 8'hFF;
            13'd4103: data <= 8'hF0;
            13'd4104: data <= 8'h00;
            13'd4105: data <= 8'h00;
            13'd4106: data <= 8'h00;
            13'd4107: data <= 8'h00;
            13'd4108: data <= 8'h00;
            13'd4109: data <= 8'h00;
            13'd4110: data <= 8'h00;
            13'd4111: data <= 8'h00;
            13'd4112: data <= 8'h00;
            13'd4113: data <= 8'h00;
            13'd4114: data <= 8'h00;
            13'd4115: data <= 8'h03;
            13'd4116: data <= 8'hFF;
            13'd4117: data <= 8'hFF;
            13'd4118: data <= 8'hFF;
            13'd4119: data <= 8'hF0;
            13'd4120: data <= 8'h7F;
            13'd4121: data <= 8'hFF;
            13'd4122: data <= 8'hFF;
            13'd4123: data <= 8'hFF;
            13'd4124: data <= 8'hFF;
            13'd4125: data <= 8'hFF;
            13'd4126: data <= 8'hFF;
            13'd4127: data <= 8'hFF;
            13'd4128: data <= 8'hFF;
            13'd4129: data <= 8'hFF;
            13'd4130: data <= 8'hFF;
            13'd4131: data <= 8'hFF;
            13'd4132: data <= 8'hFF;
            13'd4133: data <= 8'hF0;
            13'd4134: data <= 8'h00;
            13'd4135: data <= 8'h00;
            13'd4136: data <= 8'h00;
            13'd4137: data <= 8'h00;
            13'd4138: data <= 8'h00;
            13'd4139: data <= 8'h00;
            13'd4140: data <= 8'h00;
            13'd4141: data <= 8'h00;
            13'd4142: data <= 8'h00;
            13'd4143: data <= 8'h00;
            13'd4144: data <= 8'h00;
            13'd4145: data <= 8'h03;
            13'd4146: data <= 8'hFF;
            13'd4147: data <= 8'hFF;
            13'd4148: data <= 8'hFF;
            13'd4149: data <= 8'hF0;
            13'd4150: data <= 8'h7F;
            13'd4151: data <= 8'hFF;
            13'd4152: data <= 8'hFF;
            13'd4153: data <= 8'hFF;
            13'd4154: data <= 8'hFF;
            13'd4155: data <= 8'hFF;
            13'd4156: data <= 8'hFF;
            13'd4157: data <= 8'hFF;
            13'd4158: data <= 8'hFF;
            13'd4159: data <= 8'hFF;
            13'd4160: data <= 8'hFF;
            13'd4161: data <= 8'hFF;
            13'd4162: data <= 8'hFF;
            13'd4163: data <= 8'hF0;
            13'd4164: data <= 8'h00;
            13'd4165: data <= 8'h00;
            13'd4166: data <= 8'h00;
            13'd4167: data <= 8'h00;
            13'd4168: data <= 8'h00;
            13'd4169: data <= 8'h00;
            13'd4170: data <= 8'h00;
            13'd4171: data <= 8'h00;
            13'd4172: data <= 8'h00;
            13'd4173: data <= 8'h00;
            13'd4174: data <= 8'h00;
            13'd4175: data <= 8'h03;
            13'd4176: data <= 8'hFF;
            13'd4177: data <= 8'hFF;
            13'd4178: data <= 8'hFF;
            13'd4179: data <= 8'hF0;
            13'd4180: data <= 8'h7F;
            13'd4181: data <= 8'hFF;
            13'd4182: data <= 8'hFF;
            13'd4183: data <= 8'hFF;
            13'd4184: data <= 8'hFF;
            13'd4185: data <= 8'hFF;
            13'd4186: data <= 8'hFF;
            13'd4187: data <= 8'hFF;
            13'd4188: data <= 8'hFF;
            13'd4189: data <= 8'hFF;
            13'd4190: data <= 8'hFF;
            13'd4191: data <= 8'hFF;
            13'd4192: data <= 8'hFF;
            13'd4193: data <= 8'hF0;
            13'd4194: data <= 8'h00;
            13'd4195: data <= 8'h00;
            13'd4196: data <= 8'h00;
            13'd4197: data <= 8'h00;
            13'd4198: data <= 8'h00;
            13'd4199: data <= 8'h00;
            13'd4200: data <= 8'h00;
            13'd4201: data <= 8'h00;
            13'd4202: data <= 8'h00;
            13'd4203: data <= 8'h00;
            13'd4204: data <= 8'h00;
            13'd4205: data <= 8'h03;
            13'd4206: data <= 8'hFF;
            13'd4207: data <= 8'hFF;
            13'd4208: data <= 8'hFF;
            13'd4209: data <= 8'hF0;
            13'd4210: data <= 8'h7F;
            13'd4211: data <= 8'hFF;
            13'd4212: data <= 8'hFF;
            13'd4213: data <= 8'hFF;
            13'd4214: data <= 8'hFF;
            13'd4215: data <= 8'hFF;
            13'd4216: data <= 8'hFF;
            13'd4217: data <= 8'hFF;
            13'd4218: data <= 8'hFF;
            13'd4219: data <= 8'hFF;
            13'd4220: data <= 8'hFF;
            13'd4221: data <= 8'hFF;
            13'd4222: data <= 8'hFF;
            13'd4223: data <= 8'hF0;
            13'd4224: data <= 8'h00;
            13'd4225: data <= 8'h00;
            13'd4226: data <= 8'h00;
            13'd4227: data <= 8'h00;
            13'd4228: data <= 8'h00;
            13'd4229: data <= 8'h00;
            13'd4230: data <= 8'h00;
            13'd4231: data <= 8'h00;
            13'd4232: data <= 8'h00;
            13'd4233: data <= 8'h00;
            13'd4234: data <= 8'h00;
            13'd4235: data <= 8'h03;
            13'd4236: data <= 8'hFF;
            13'd4237: data <= 8'hFF;
            13'd4238: data <= 8'hFF;
            13'd4239: data <= 8'hF0;
            13'd4240: data <= 8'h7F;
            13'd4241: data <= 8'hFF;
            13'd4242: data <= 8'hFF;
            13'd4243: data <= 8'hFF;
            13'd4244: data <= 8'hFF;
            13'd4245: data <= 8'hFF;
            13'd4246: data <= 8'hFF;
            13'd4247: data <= 8'hFF;
            13'd4248: data <= 8'hFF;
            13'd4249: data <= 8'hFF;
            13'd4250: data <= 8'hFF;
            13'd4251: data <= 8'hFF;
            13'd4252: data <= 8'hFF;
            13'd4253: data <= 8'hF0;
            13'd4254: data <= 8'h00;
            13'd4255: data <= 8'h00;
            13'd4256: data <= 8'h00;
            13'd4257: data <= 8'h00;
            13'd4258: data <= 8'h00;
            13'd4259: data <= 8'h00;
            13'd4260: data <= 8'h00;
            13'd4261: data <= 8'h00;
            13'd4262: data <= 8'h00;
            13'd4263: data <= 8'h00;
            13'd4264: data <= 8'h00;
            13'd4265: data <= 8'h03;
            13'd4266: data <= 8'hFF;
            13'd4267: data <= 8'hFF;
            13'd4268: data <= 8'hFF;
            13'd4269: data <= 8'hF0;
            13'd4270: data <= 8'h7F;
            13'd4271: data <= 8'hFF;
            13'd4272: data <= 8'hFF;
            13'd4273: data <= 8'hFF;
            13'd4274: data <= 8'hFF;
            13'd4275: data <= 8'hFF;
            13'd4276: data <= 8'hFF;
            13'd4277: data <= 8'hFF;
            13'd4278: data <= 8'hFF;
            13'd4279: data <= 8'hFF;
            13'd4280: data <= 8'hFF;
            13'd4281: data <= 8'hFF;
            13'd4282: data <= 8'hFF;
            13'd4283: data <= 8'hF8;
            13'd4284: data <= 8'h00;
            13'd4285: data <= 8'h00;
            13'd4286: data <= 8'h00;
            13'd4287: data <= 8'h00;
            13'd4288: data <= 8'h00;
            13'd4289: data <= 8'h00;
            13'd4290: data <= 8'h00;
            13'd4291: data <= 8'h00;
            13'd4292: data <= 8'h00;
            13'd4293: data <= 8'h00;
            13'd4294: data <= 8'h00;
            13'd4295: data <= 8'h03;
            13'd4296: data <= 8'hFF;
            13'd4297: data <= 8'hFF;
            13'd4298: data <= 8'hFF;
            13'd4299: data <= 8'hE0;
            13'd4300: data <= 8'h7F;
            13'd4301: data <= 8'hFF;
            13'd4302: data <= 8'hFF;
            13'd4303: data <= 8'hFF;
            13'd4304: data <= 8'hFF;
            13'd4305: data <= 8'hFF;
            13'd4306: data <= 8'hFF;
            13'd4307: data <= 8'hFF;
            13'd4308: data <= 8'hFF;
            13'd4309: data <= 8'hFF;
            13'd4310: data <= 8'hFF;
            13'd4311: data <= 8'hFF;
            13'd4312: data <= 8'hFF;
            13'd4313: data <= 8'hF8;
            13'd4314: data <= 8'h00;
            13'd4315: data <= 8'h00;
            13'd4316: data <= 8'h00;
            13'd4317: data <= 8'h00;
            13'd4318: data <= 8'h00;
            13'd4319: data <= 8'h00;
            13'd4320: data <= 8'h00;
            13'd4321: data <= 8'h00;
            13'd4322: data <= 8'h00;
            13'd4323: data <= 8'h00;
            13'd4324: data <= 8'h00;
            13'd4325: data <= 8'h03;
            13'd4326: data <= 8'hFF;
            13'd4327: data <= 8'hFF;
            13'd4328: data <= 8'hFF;
            13'd4329: data <= 8'hE0;
            13'd4330: data <= 8'h7F;
            13'd4331: data <= 8'hFF;
            13'd4332: data <= 8'hFF;
            13'd4333: data <= 8'hFF;
            13'd4334: data <= 8'hFF;
            13'd4335: data <= 8'hFF;
            13'd4336: data <= 8'hFF;
            13'd4337: data <= 8'hFF;
            13'd4338: data <= 8'hFF;
            13'd4339: data <= 8'hFF;
            13'd4340: data <= 8'hFF;
            13'd4341: data <= 8'hFF;
            13'd4342: data <= 8'hFF;
            13'd4343: data <= 8'hF8;
            13'd4344: data <= 8'h00;
            13'd4345: data <= 8'h00;
            13'd4346: data <= 8'h00;
            13'd4347: data <= 8'h00;
            13'd4348: data <= 8'h00;
            13'd4349: data <= 8'h00;
            13'd4350: data <= 8'h00;
            13'd4351: data <= 8'h00;
            13'd4352: data <= 8'h00;
            13'd4353: data <= 8'h00;
            13'd4354: data <= 8'h00;
            13'd4355: data <= 8'h03;
            13'd4356: data <= 8'hFF;
            13'd4357: data <= 8'hFF;
            13'd4358: data <= 8'hFF;
            13'd4359: data <= 8'hE0;
            13'd4360: data <= 8'h7F;
            13'd4361: data <= 8'hFF;
            13'd4362: data <= 8'hFF;
            13'd4363: data <= 8'hFF;
            13'd4364: data <= 8'hFF;
            13'd4365: data <= 8'hFF;
            13'd4366: data <= 8'hFF;
            13'd4367: data <= 8'hFF;
            13'd4368: data <= 8'hFF;
            13'd4369: data <= 8'hFF;
            13'd4370: data <= 8'hFF;
            13'd4371: data <= 8'hFF;
            13'd4372: data <= 8'hFF;
            13'd4373: data <= 8'hF8;
            13'd4374: data <= 8'h00;
            13'd4375: data <= 8'h00;
            13'd4376: data <= 8'h00;
            13'd4377: data <= 8'h00;
            13'd4378: data <= 8'h00;
            13'd4379: data <= 8'h00;
            13'd4380: data <= 8'h00;
            13'd4381: data <= 8'h00;
            13'd4382: data <= 8'h00;
            13'd4383: data <= 8'h00;
            13'd4384: data <= 8'h00;
            13'd4385: data <= 8'h03;
            13'd4386: data <= 8'hFF;
            13'd4387: data <= 8'hFF;
            13'd4388: data <= 8'hFF;
            13'd4389: data <= 8'hE0;
            13'd4390: data <= 8'h7F;
            13'd4391: data <= 8'hFF;
            13'd4392: data <= 8'hFF;
            13'd4393: data <= 8'hFF;
            13'd4394: data <= 8'hFF;
            13'd4395: data <= 8'hFF;
            13'd4396: data <= 8'hFF;
            13'd4397: data <= 8'hFF;
            13'd4398: data <= 8'hFF;
            13'd4399: data <= 8'hFF;
            13'd4400: data <= 8'hFF;
            13'd4401: data <= 8'hFF;
            13'd4402: data <= 8'hFF;
            13'd4403: data <= 8'hF8;
            13'd4404: data <= 8'h00;
            13'd4405: data <= 8'h00;
            13'd4406: data <= 8'h00;
            13'd4407: data <= 8'h00;
            13'd4408: data <= 8'h00;
            13'd4409: data <= 8'h00;
            13'd4410: data <= 8'h00;
            13'd4411: data <= 8'h00;
            13'd4412: data <= 8'h00;
            13'd4413: data <= 8'h00;
            13'd4414: data <= 8'h00;
            13'd4415: data <= 8'h03;
            13'd4416: data <= 8'hFF;
            13'd4417: data <= 8'hFF;
            13'd4418: data <= 8'hFF;
            13'd4419: data <= 8'hF0;
            13'd4420: data <= 8'hFF;
            13'd4421: data <= 8'hFF;
            13'd4422: data <= 8'hFF;
            13'd4423: data <= 8'hFF;
            13'd4424: data <= 8'hFF;
            13'd4425: data <= 8'hFF;
            13'd4426: data <= 8'hFF;
            13'd4427: data <= 8'hFF;
            13'd4428: data <= 8'hFF;
            13'd4429: data <= 8'hFF;
            13'd4430: data <= 8'hFF;
            13'd4431: data <= 8'hFF;
            13'd4432: data <= 8'hFF;
            13'd4433: data <= 8'hFC;
            13'd4434: data <= 8'h00;
            13'd4435: data <= 8'h00;
            13'd4436: data <= 8'h00;
            13'd4437: data <= 8'h00;
            13'd4438: data <= 8'h00;
            13'd4439: data <= 8'h00;
            13'd4440: data <= 8'h00;
            13'd4441: data <= 8'h00;
            13'd4442: data <= 8'h00;
            13'd4443: data <= 8'h00;
            13'd4444: data <= 8'h00;
            13'd4445: data <= 8'h03;
            13'd4446: data <= 8'hFF;
            13'd4447: data <= 8'hFF;
            13'd4448: data <= 8'hFF;
            13'd4449: data <= 8'hFF;
            13'd4450: data <= 8'hFF;
            13'd4451: data <= 8'hFF;
            13'd4452: data <= 8'hFF;
            13'd4453: data <= 8'hFF;
            13'd4454: data <= 8'hFF;
            13'd4455: data <= 8'hFF;
            13'd4456: data <= 8'hFF;
            13'd4457: data <= 8'hFF;
            13'd4458: data <= 8'hFF;
            13'd4459: data <= 8'hFF;
            13'd4460: data <= 8'hFF;
            13'd4461: data <= 8'hFF;
            13'd4462: data <= 8'hFF;
            13'd4463: data <= 8'hFF;
            13'd4464: data <= 8'h80;
            13'd4465: data <= 8'h00;
            13'd4466: data <= 8'h00;
            13'd4467: data <= 8'h00;
            13'd4468: data <= 8'h00;
            13'd4469: data <= 8'h00;
            13'd4470: data <= 8'h00;
            13'd4471: data <= 8'h00;
            13'd4472: data <= 8'h00;
            13'd4473: data <= 8'h00;
            13'd4474: data <= 8'h00;
            13'd4475: data <= 8'h03;
            13'd4476: data <= 8'hFF;
            13'd4477: data <= 8'hFF;
            13'd4478: data <= 8'hFF;
            13'd4479: data <= 8'hFF;
            13'd4480: data <= 8'hFF;
            13'd4481: data <= 8'hFF;
            13'd4482: data <= 8'hFF;
            13'd4483: data <= 8'hFF;
            13'd4484: data <= 8'hFF;
            13'd4485: data <= 8'hFF;
            13'd4486: data <= 8'hFF;
            13'd4487: data <= 8'hFF;
            13'd4488: data <= 8'hFF;
            13'd4489: data <= 8'hFF;
            13'd4490: data <= 8'hFF;
            13'd4491: data <= 8'hFF;
            13'd4492: data <= 8'hFF;
            13'd4493: data <= 8'hFF;
            13'd4494: data <= 8'h80;
            13'd4495: data <= 8'h00;
            13'd4496: data <= 8'h00;
            13'd4497: data <= 8'h00;
            13'd4498: data <= 8'h00;
            13'd4499: data <= 8'h00;
            13'd4500: data <= 8'h00;
            13'd4501: data <= 8'h00;
            13'd4502: data <= 8'h00;
            13'd4503: data <= 8'h00;
            13'd4504: data <= 8'h00;
            13'd4505: data <= 8'h03;
            13'd4506: data <= 8'hFF;
            13'd4507: data <= 8'hFF;
            13'd4508: data <= 8'hFF;
            13'd4509: data <= 8'hFF;
            13'd4510: data <= 8'hFF;
            13'd4511: data <= 8'hFF;
            13'd4512: data <= 8'hFF;
            13'd4513: data <= 8'hFF;
            13'd4514: data <= 8'hFF;
            13'd4515: data <= 8'hFF;
            13'd4516: data <= 8'hFF;
            13'd4517: data <= 8'hFF;
            13'd4518: data <= 8'hFF;
            13'd4519: data <= 8'hFF;
            13'd4520: data <= 8'hFF;
            13'd4521: data <= 8'hFF;
            13'd4522: data <= 8'hFF;
            13'd4523: data <= 8'hFF;
            13'd4524: data <= 8'h80;
            13'd4525: data <= 8'h00;
            13'd4526: data <= 8'h00;
            13'd4527: data <= 8'h00;
            13'd4528: data <= 8'h00;
            13'd4529: data <= 8'h00;
            13'd4530: data <= 8'h00;
            13'd4531: data <= 8'h00;
            13'd4532: data <= 8'h00;
            13'd4533: data <= 8'h00;
            13'd4534: data <= 8'h00;
            13'd4535: data <= 8'h03;
            13'd4536: data <= 8'hFF;
            13'd4537: data <= 8'hFF;
            13'd4538: data <= 8'hFF;
            13'd4539: data <= 8'hFF;
            13'd4540: data <= 8'hFF;
            13'd4541: data <= 8'hFF;
            13'd4542: data <= 8'hFF;
            13'd4543: data <= 8'hFF;
            13'd4544: data <= 8'hFF;
            13'd4545: data <= 8'hFF;
            13'd4546: data <= 8'hFF;
            13'd4547: data <= 8'hFF;
            13'd4548: data <= 8'hFF;
            13'd4549: data <= 8'hFF;
            13'd4550: data <= 8'hFF;
            13'd4551: data <= 8'hFF;
            13'd4552: data <= 8'hFF;
            13'd4553: data <= 8'hFF;
            13'd4554: data <= 8'h80;
            13'd4555: data <= 8'h00;
            13'd4556: data <= 8'h00;
            13'd4557: data <= 8'h00;
            13'd4558: data <= 8'h00;
            13'd4559: data <= 8'h00;
            13'd4560: data <= 8'h00;
            13'd4561: data <= 8'h00;
            13'd4562: data <= 8'h00;
            13'd4563: data <= 8'h00;
            13'd4564: data <= 8'h00;
            13'd4565: data <= 8'h03;
            13'd4566: data <= 8'hFF;
            13'd4567: data <= 8'hFF;
            13'd4568: data <= 8'hFF;
            13'd4569: data <= 8'hFF;
            13'd4570: data <= 8'hFF;
            13'd4571: data <= 8'hFF;
            13'd4572: data <= 8'hFF;
            13'd4573: data <= 8'hFF;
            13'd4574: data <= 8'hFF;
            13'd4575: data <= 8'hFF;
            13'd4576: data <= 8'hFF;
            13'd4577: data <= 8'hFF;
            13'd4578: data <= 8'hFF;
            13'd4579: data <= 8'hFF;
            13'd4580: data <= 8'hFF;
            13'd4581: data <= 8'hFF;
            13'd4582: data <= 8'hFF;
            13'd4583: data <= 8'hFF;
            13'd4584: data <= 8'h80;
            13'd4585: data <= 8'h00;
            13'd4586: data <= 8'h00;
            13'd4587: data <= 8'h00;
            13'd4588: data <= 8'h00;
            13'd4589: data <= 8'h00;
            13'd4590: data <= 8'h00;
            13'd4591: data <= 8'h00;
            13'd4592: data <= 8'h00;
            13'd4593: data <= 8'h00;
            13'd4594: data <= 8'h00;
            13'd4595: data <= 8'h03;
            13'd4596: data <= 8'hFF;
            13'd4597: data <= 8'hFF;
            13'd4598: data <= 8'hFF;
            13'd4599: data <= 8'hFF;
            13'd4600: data <= 8'hFF;
            13'd4601: data <= 8'hFF;
            13'd4602: data <= 8'hFF;
            13'd4603: data <= 8'hFF;
            13'd4604: data <= 8'hFF;
            13'd4605: data <= 8'hFF;
            13'd4606: data <= 8'hFF;
            13'd4607: data <= 8'hFF;
            13'd4608: data <= 8'hFF;
            13'd4609: data <= 8'hFF;
            13'd4610: data <= 8'hFF;
            13'd4611: data <= 8'hFF;
            13'd4612: data <= 8'hFF;
            13'd4613: data <= 8'hFF;
            13'd4614: data <= 8'h80;
            13'd4615: data <= 8'h00;
            13'd4616: data <= 8'h00;
            13'd4617: data <= 8'h00;
            13'd4618: data <= 8'h00;
            13'd4619: data <= 8'h00;
            13'd4620: data <= 8'h00;
            13'd4621: data <= 8'h00;
            13'd4622: data <= 8'h00;
            13'd4623: data <= 8'h00;
            13'd4624: data <= 8'h00;
            13'd4625: data <= 8'h03;
            13'd4626: data <= 8'hFF;
            13'd4627: data <= 8'hFF;
            13'd4628: data <= 8'hFF;
            13'd4629: data <= 8'hFF;
            13'd4630: data <= 8'hFF;
            13'd4631: data <= 8'hFF;
            13'd4632: data <= 8'hFF;
            13'd4633: data <= 8'hFF;
            13'd4634: data <= 8'hFF;
            13'd4635: data <= 8'hFF;
            13'd4636: data <= 8'hFF;
            13'd4637: data <= 8'hFF;
            13'd4638: data <= 8'hFF;
            13'd4639: data <= 8'hFF;
            13'd4640: data <= 8'hFF;
            13'd4641: data <= 8'hFF;
            13'd4642: data <= 8'hFF;
            13'd4643: data <= 8'hFF;
            13'd4644: data <= 8'h80;
            13'd4645: data <= 8'h00;
            13'd4646: data <= 8'h00;
            13'd4647: data <= 8'h00;
            13'd4648: data <= 8'h00;
            13'd4649: data <= 8'h00;
            13'd4650: data <= 8'h00;
            13'd4651: data <= 8'h00;
            13'd4652: data <= 8'h00;
            13'd4653: data <= 8'h00;
            13'd4654: data <= 8'h00;
            13'd4655: data <= 8'h03;
            13'd4656: data <= 8'hFF;
            13'd4657: data <= 8'hFF;
            13'd4658: data <= 8'hFF;
            13'd4659: data <= 8'hFF;
            13'd4660: data <= 8'hFF;
            13'd4661: data <= 8'hFF;
            13'd4662: data <= 8'hFF;
            13'd4663: data <= 8'hFF;
            13'd4664: data <= 8'hFF;
            13'd4665: data <= 8'hFF;
            13'd4666: data <= 8'hFF;
            13'd4667: data <= 8'hFF;
            13'd4668: data <= 8'h8F;
            13'd4669: data <= 8'hFF;
            13'd4670: data <= 8'hFF;
            13'd4671: data <= 8'hFF;
            13'd4672: data <= 8'hFF;
            13'd4673: data <= 8'hFF;
            13'd4674: data <= 8'h80;
            13'd4675: data <= 8'h00;
            13'd4676: data <= 8'h00;
            13'd4677: data <= 8'h00;
            13'd4678: data <= 8'h00;
            13'd4679: data <= 8'h00;
            13'd4680: data <= 8'h00;
            13'd4681: data <= 8'h00;
            13'd4682: data <= 8'h00;
            13'd4683: data <= 8'h00;
            13'd4684: data <= 8'h00;
            13'd4685: data <= 8'h03;
            13'd4686: data <= 8'hFF;
            13'd4687: data <= 8'hFF;
            13'd4688: data <= 8'hFF;
            13'd4689: data <= 8'hFF;
            13'd4690: data <= 8'hFB;
            13'd4691: data <= 8'hFF;
            13'd4692: data <= 8'hFF;
            13'd4693: data <= 8'hFF;
            13'd4694: data <= 8'hFE;
            13'd4695: data <= 8'hFF;
            13'd4696: data <= 8'hFF;
            13'd4697: data <= 8'hF8;
            13'd4698: data <= 8'h07;
            13'd4699: data <= 8'hFF;
            13'd4700: data <= 8'hFF;
            13'd4701: data <= 8'hFF;
            13'd4702: data <= 8'hFF;
            13'd4703: data <= 8'hFF;
            13'd4704: data <= 8'h80;
            13'd4705: data <= 8'h00;
            13'd4706: data <= 8'h00;
            13'd4707: data <= 8'h00;
            13'd4708: data <= 8'h00;
            13'd4709: data <= 8'h00;
            13'd4710: data <= 8'h00;
            13'd4711: data <= 8'h00;
            13'd4712: data <= 8'h00;
            13'd4713: data <= 8'h00;
            13'd4714: data <= 8'h00;
            13'd4715: data <= 8'h03;
            13'd4716: data <= 8'hFF;
            13'd4717: data <= 8'hE0;
            13'd4718: data <= 8'h00;
            13'd4719: data <= 8'h3C;
            13'd4720: data <= 8'h0B;
            13'd4721: data <= 8'h7F;
            13'd4722: data <= 8'hFF;
            13'd4723: data <= 8'hFF;
            13'd4724: data <= 8'hFC;
            13'd4725: data <= 8'h7F;
            13'd4726: data <= 8'hFF;
            13'd4727: data <= 8'hC3;
            13'd4728: data <= 8'hF1;
            13'd4729: data <= 8'hFF;
            13'd4730: data <= 8'hFF;
            13'd4731: data <= 8'hE0;
            13'd4732: data <= 8'h1F;
            13'd4733: data <= 8'hFF;
            13'd4734: data <= 8'h80;
            13'd4735: data <= 8'h00;
            13'd4736: data <= 8'h00;
            13'd4737: data <= 8'h00;
            13'd4738: data <= 8'h00;
            13'd4739: data <= 8'h00;
            13'd4740: data <= 8'h00;
            13'd4741: data <= 8'h00;
            13'd4742: data <= 8'h00;
            13'd4743: data <= 8'h00;
            13'd4744: data <= 8'h00;
            13'd4745: data <= 8'h03;
            13'd4746: data <= 8'hFF;
            13'd4747: data <= 8'hFF;
            13'd4748: data <= 8'h77;
            13'd4749: data <= 8'hF0;
            13'd4750: data <= 8'h7B;
            13'd4751: data <= 8'h1F;
            13'd4752: data <= 8'hFF;
            13'd4753: data <= 8'hFE;
            13'd4754: data <= 8'h00;
            13'd4755: data <= 8'h00;
            13'd4756: data <= 8'hFF;
            13'd4757: data <= 8'h9F;
            13'd4758: data <= 8'hFC;
            13'd4759: data <= 8'h3F;
            13'd4760: data <= 8'hF8;
            13'd4761: data <= 8'h7F;
            13'd4762: data <= 8'h9F;
            13'd4763: data <= 8'hFF;
            13'd4764: data <= 8'h80;
            13'd4765: data <= 8'h00;
            13'd4766: data <= 8'h00;
            13'd4767: data <= 8'h00;
            13'd4768: data <= 8'h00;
            13'd4769: data <= 8'h00;
            13'd4770: data <= 8'h00;
            13'd4771: data <= 8'h00;
            13'd4772: data <= 8'h00;
            13'd4773: data <= 8'h00;
            13'd4774: data <= 8'h00;
            13'd4775: data <= 8'h03;
            13'd4776: data <= 8'hFF;
            13'd4777: data <= 8'hFF;
            13'd4778: data <= 8'h77;
            13'd4779: data <= 8'hFE;
            13'd4780: data <= 8'h7B;
            13'd4781: data <= 8'hDF;
            13'd4782: data <= 8'hFF;
            13'd4783: data <= 8'hFF;
            13'd4784: data <= 8'hFE;
            13'd4785: data <= 8'hFF;
            13'd4786: data <= 8'hFF;
            13'd4787: data <= 8'h3F;
            13'd4788: data <= 8'hFF;
            13'd4789: data <= 8'h9F;
            13'd4790: data <= 8'hFB;
            13'd4791: data <= 8'h37;
            13'd4792: data <= 8'h9F;
            13'd4793: data <= 8'hFF;
            13'd4794: data <= 8'h80;
            13'd4795: data <= 8'h00;
            13'd4796: data <= 8'h00;
            13'd4797: data <= 8'h00;
            13'd4798: data <= 8'h00;
            13'd4799: data <= 8'h00;
            13'd4800: data <= 8'h00;
            13'd4801: data <= 8'h00;
            13'd4802: data <= 8'h00;
            13'd4803: data <= 8'h00;
            13'd4804: data <= 8'h00;
            13'd4805: data <= 8'h03;
            13'd4806: data <= 8'hFF;
            13'd4807: data <= 8'hF0;
            13'd4808: data <= 8'h00;
            13'd4809: data <= 8'h3E;
            13'd4810: data <= 8'h7B;
            13'd4811: data <= 8'hFF;
            13'd4812: data <= 8'hFF;
            13'd4813: data <= 8'hFF;
            13'd4814: data <= 8'hC0;
            13'd4815: data <= 8'h0F;
            13'd4816: data <= 8'hFE;
            13'd4817: data <= 8'h7F;
            13'd4818: data <= 8'hFF;
            13'd4819: data <= 8'h9F;
            13'd4820: data <= 8'hFB;
            13'd4821: data <= 8'h37;
            13'd4822: data <= 8'h9F;
            13'd4823: data <= 8'hFF;
            13'd4824: data <= 8'h80;
            13'd4825: data <= 8'h00;
            13'd4826: data <= 8'h00;
            13'd4827: data <= 8'h00;
            13'd4828: data <= 8'h00;
            13'd4829: data <= 8'h00;
            13'd4830: data <= 8'h00;
            13'd4831: data <= 8'h00;
            13'd4832: data <= 8'h00;
            13'd4833: data <= 8'h00;
            13'd4834: data <= 8'h00;
            13'd4835: data <= 8'h03;
            13'd4836: data <= 8'hFF;
            13'd4837: data <= 8'hE7;
            13'd4838: data <= 8'h77;
            13'd4839: data <= 8'h30;
            13'd4840: data <= 8'h00;
            13'd4841: data <= 8'h0F;
            13'd4842: data <= 8'hFF;
            13'd4843: data <= 8'hFF;
            13'd4844: data <= 8'h80;
            13'd4845: data <= 8'h03;
            13'd4846: data <= 8'hFE;
            13'd4847: data <= 8'hEF;
            13'd4848: data <= 8'hFF;
            13'd4849: data <= 8'hDF;
            13'd4850: data <= 8'hFB;
            13'd4851: data <= 8'h27;
            13'd4852: data <= 8'h9F;
            13'd4853: data <= 8'hFF;
            13'd4854: data <= 8'h80;
            13'd4855: data <= 8'h00;
            13'd4856: data <= 8'h00;
            13'd4857: data <= 8'h00;
            13'd4858: data <= 8'h00;
            13'd4859: data <= 8'h00;
            13'd4860: data <= 8'h00;
            13'd4861: data <= 8'h00;
            13'd4862: data <= 8'h00;
            13'd4863: data <= 8'h00;
            13'd4864: data <= 8'h00;
            13'd4865: data <= 8'h03;
            13'd4866: data <= 8'hFF;
            13'd4867: data <= 8'hE7;
            13'd4868: data <= 8'h77;
            13'd4869: data <= 8'h30;
            13'd4870: data <= 8'h00;
            13'd4871: data <= 8'h07;
            13'd4872: data <= 8'hFF;
            13'd4873: data <= 8'hFF;
            13'd4874: data <= 8'h9F;
            13'd4875: data <= 8'hF3;
            13'd4876: data <= 8'hFE;
            13'd4877: data <= 8'hFF;
            13'd4878: data <= 8'hFF;
            13'd4879: data <= 8'hCF;
            13'd4880: data <= 8'hFB;
            13'd4881: data <= 8'h27;
            13'd4882: data <= 8'hBF;
            13'd4883: data <= 8'hFF;
            13'd4884: data <= 8'h80;
            13'd4885: data <= 8'h00;
            13'd4886: data <= 8'h00;
            13'd4887: data <= 8'h00;
            13'd4888: data <= 8'h00;
            13'd4889: data <= 8'h00;
            13'd4890: data <= 8'h00;
            13'd4891: data <= 8'h00;
            13'd4892: data <= 8'h00;
            13'd4893: data <= 8'h00;
            13'd4894: data <= 8'h00;
            13'd4895: data <= 8'h03;
            13'd4896: data <= 8'hFF;
            13'd4897: data <= 8'hE0;
            13'd4898: data <= 8'h00;
            13'd4899: data <= 8'h3E;
            13'd4900: data <= 8'h79;
            13'd4901: data <= 8'hFC;
            13'd4902: data <= 8'h00;
            13'd4903: data <= 8'h03;
            13'd4904: data <= 8'h80;
            13'd4905: data <= 8'h03;
            13'd4906: data <= 8'hFE;
            13'd4907: data <= 8'hFF;
            13'd4908: data <= 8'hFF;
            13'd4909: data <= 8'hE7;
            13'd4910: data <= 8'hFB;
            13'd4911: data <= 8'h27;
            13'd4912: data <= 8'hBF;
            13'd4913: data <= 8'hFF;
            13'd4914: data <= 8'h80;
            13'd4915: data <= 8'h00;
            13'd4916: data <= 8'h00;
            13'd4917: data <= 8'h00;
            13'd4918: data <= 8'h00;
            13'd4919: data <= 8'h00;
            13'd4920: data <= 8'h00;
            13'd4921: data <= 8'h00;
            13'd4922: data <= 8'h00;
            13'd4923: data <= 8'h00;
            13'd4924: data <= 8'h00;
            13'd4925: data <= 8'h03;
            13'd4926: data <= 8'hFF;
            13'd4927: data <= 8'hF7;
            13'd4928: data <= 8'h7F;
            13'd4929: data <= 8'h3E;
            13'd4930: data <= 8'h79;
            13'd4931: data <= 8'hC8;
            13'd4932: data <= 8'h00;
            13'd4933: data <= 8'h03;
            13'd4934: data <= 8'h9F;
            13'd4935: data <= 8'hF3;
            13'd4936: data <= 8'hFE;
            13'd4937: data <= 8'hE3;
            13'd4938: data <= 8'hFF;
            13'd4939: data <= 8'hF7;
            13'd4940: data <= 8'hFB;
            13'd4941: data <= 8'h20;
            13'd4942: data <= 8'h0F;
            13'd4943: data <= 8'hFF;
            13'd4944: data <= 8'h80;
            13'd4945: data <= 8'h00;
            13'd4946: data <= 8'h00;
            13'd4947: data <= 8'h00;
            13'd4948: data <= 8'h00;
            13'd4949: data <= 8'h00;
            13'd4950: data <= 8'h00;
            13'd4951: data <= 8'h00;
            13'd4952: data <= 8'h00;
            13'd4953: data <= 8'h00;
            13'd4954: data <= 8'h00;
            13'd4955: data <= 8'h03;
            13'd4956: data <= 8'hFF;
            13'd4957: data <= 8'hFF;
            13'd4958: data <= 8'h7F;
            13'd4959: data <= 8'hFE;
            13'd4960: data <= 8'h0D;
            13'd4961: data <= 8'h9F;
            13'd4962: data <= 8'hFF;
            13'd4963: data <= 8'hFF;
            13'd4964: data <= 8'h9F;
            13'd4965: data <= 8'hF3;
            13'd4966: data <= 8'hFE;
            13'd4967: data <= 8'h05;
            13'd4968: data <= 8'hFF;
            13'd4969: data <= 8'hF3;
            13'd4970: data <= 8'hFB;
            13'd4971: data <= 8'h3F;
            13'd4972: data <= 8'hEF;
            13'd4973: data <= 8'hFF;
            13'd4974: data <= 8'h80;
            13'd4975: data <= 8'h00;
            13'd4976: data <= 8'h00;
            13'd4977: data <= 8'h00;
            13'd4978: data <= 8'h00;
            13'd4979: data <= 8'h00;
            13'd4980: data <= 8'h00;
            13'd4981: data <= 8'h00;
            13'd4982: data <= 8'h00;
            13'd4983: data <= 8'h00;
            13'd4984: data <= 8'h00;
            13'd4985: data <= 8'h03;
            13'd4986: data <= 8'hFF;
            13'd4987: data <= 8'hC0;
            13'd4988: data <= 8'h00;
            13'd4989: data <= 8'h10;
            13'd4990: data <= 8'h1D;
            13'd4991: data <= 8'h3F;
            13'd4992: data <= 8'hFF;
            13'd4993: data <= 8'hFF;
            13'd4994: data <= 8'h80;
            13'd4995: data <= 8'h03;
            13'd4996: data <= 8'hFF;
            13'd4997: data <= 8'h01;
            13'd4998: data <= 8'hFF;
            13'd4999: data <= 8'hFB;
            13'd5000: data <= 8'hFB;
            13'd5001: data <= 8'h3F;
            13'd5002: data <= 8'hEF;
            13'd5003: data <= 8'hFF;
            13'd5004: data <= 8'h80;
            13'd5005: data <= 8'h00;
            13'd5006: data <= 8'h00;
            13'd5007: data <= 8'h00;
            13'd5008: data <= 8'h00;
            13'd5009: data <= 8'h00;
            13'd5010: data <= 8'h00;
            13'd5011: data <= 8'h00;
            13'd5012: data <= 8'h00;
            13'd5013: data <= 8'h00;
            13'd5014: data <= 8'h00;
            13'd5015: data <= 8'h03;
            13'd5016: data <= 8'hFF;
            13'd5017: data <= 8'hFC;
            13'd5018: data <= 8'hF9;
            13'd5019: data <= 8'hF2;
            13'd5020: data <= 8'h7C;
            13'd5021: data <= 8'h7F;
            13'd5022: data <= 8'hFF;
            13'd5023: data <= 8'hFF;
            13'd5024: data <= 8'h9F;
            13'd5025: data <= 8'hF3;
            13'd5026: data <= 8'hFF;
            13'd5027: data <= 8'h9F;
            13'd5028: data <= 8'hFF;
            13'd5029: data <= 8'hFB;
            13'd5030: data <= 8'hFB;
            13'd5031: data <= 8'h3F;
            13'd5032: data <= 8'hEF;
            13'd5033: data <= 8'hFF;
            13'd5034: data <= 8'h80;
            13'd5035: data <= 8'h00;
            13'd5036: data <= 8'h00;
            13'd5037: data <= 8'h00;
            13'd5038: data <= 8'h00;
            13'd5039: data <= 8'h00;
            13'd5040: data <= 8'h00;
            13'd5041: data <= 8'h00;
            13'd5042: data <= 8'h00;
            13'd5043: data <= 8'h00;
            13'd5044: data <= 8'h00;
            13'd5045: data <= 8'h03;
            13'd5046: data <= 8'hFF;
            13'd5047: data <= 8'hFD;
            13'd5048: data <= 8'hFB;
            13'd5049: data <= 8'hFE;
            13'd5050: data <= 8'h7C;
            13'd5051: data <= 8'hFF;
            13'd5052: data <= 8'hFF;
            13'd5053: data <= 8'hFF;
            13'd5054: data <= 8'h80;
            13'd5055: data <= 8'h03;
            13'd5056: data <= 8'hFF;
            13'd5057: data <= 8'hAD;
            13'd5058: data <= 8'hFF;
            13'd5059: data <= 8'hF9;
            13'd5060: data <= 8'hF8;
            13'd5061: data <= 8'h00;
            13'd5062: data <= 8'h2F;
            13'd5063: data <= 8'hFF;
            13'd5064: data <= 8'h80;
            13'd5065: data <= 8'h00;
            13'd5066: data <= 8'h00;
            13'd5067: data <= 8'h00;
            13'd5068: data <= 8'h00;
            13'd5069: data <= 8'h00;
            13'd5070: data <= 8'h00;
            13'd5071: data <= 8'h00;
            13'd5072: data <= 8'h00;
            13'd5073: data <= 8'h00;
            13'd5074: data <= 8'h00;
            13'd5075: data <= 8'h03;
            13'd5076: data <= 8'hFF;
            13'd5077: data <= 8'hFC;
            13'd5078: data <= 8'h27;
            13'd5079: data <= 8'hFE;
            13'd5080: data <= 8'h70;
            13'd5081: data <= 8'hE7;
            13'd5082: data <= 8'hFF;
            13'd5083: data <= 8'hFF;
            13'd5084: data <= 8'h80;
            13'd5085: data <= 8'h03;
            13'd5086: data <= 8'hFF;
            13'd5087: data <= 8'hAE;
            13'd5088: data <= 8'h67;
            13'd5089: data <= 8'hFD;
            13'd5090: data <= 8'hFB;
            13'd5091: data <= 8'h3F;
            13'd5092: data <= 8'hEF;
            13'd5093: data <= 8'hFF;
            13'd5094: data <= 8'h80;
            13'd5095: data <= 8'h00;
            13'd5096: data <= 8'h00;
            13'd5097: data <= 8'h00;
            13'd5098: data <= 8'h00;
            13'd5099: data <= 8'h00;
            13'd5100: data <= 8'h00;
            13'd5101: data <= 8'h00;
            13'd5102: data <= 8'h00;
            13'd5103: data <= 8'h00;
            13'd5104: data <= 8'h00;
            13'd5105: data <= 8'h03;
            13'd5106: data <= 8'hFF;
            13'd5107: data <= 8'hFF;
            13'd5108: data <= 8'h87;
            13'd5109: data <= 8'hFE;
            13'd5110: data <= 8'h66;
            13'd5111: data <= 8'h6F;
            13'd5112: data <= 8'hFF;
            13'd5113: data <= 8'hFF;
            13'd5114: data <= 8'h9F;
            13'd5115: data <= 8'hF3;
            13'd5116: data <= 8'hFF;
            13'd5117: data <= 8'hB7;
            13'd5118: data <= 8'h8F;
            13'd5119: data <= 8'hFC;
            13'd5120: data <= 8'hFF;
            13'd5121: data <= 8'hFF;
            13'd5122: data <= 8'hEF;
            13'd5123: data <= 8'hFF;
            13'd5124: data <= 8'h80;
            13'd5125: data <= 8'h00;
            13'd5126: data <= 8'h00;
            13'd5127: data <= 8'h00;
            13'd5128: data <= 8'h00;
            13'd5129: data <= 8'h00;
            13'd5130: data <= 8'h00;
            13'd5131: data <= 8'h00;
            13'd5132: data <= 8'h00;
            13'd5133: data <= 8'h00;
            13'd5134: data <= 8'h00;
            13'd5135: data <= 8'h03;
            13'd5136: data <= 8'hFF;
            13'd5137: data <= 8'hFC;
            13'd5138: data <= 8'h30;
            13'd5139: data <= 8'h7E;
            13'd5140: data <= 8'h4F;
            13'd5141: data <= 8'h2F;
            13'd5142: data <= 8'hFF;
            13'd5143: data <= 8'hFE;
            13'd5144: data <= 8'h00;
            13'd5145: data <= 8'h00;
            13'd5146: data <= 8'hFF;
            13'd5147: data <= 8'hF7;
            13'd5148: data <= 8'hFF;
            13'd5149: data <= 8'hFC;
            13'd5150: data <= 8'hFF;
            13'd5151: data <= 8'hFC;
            13'd5152: data <= 8'h0F;
            13'd5153: data <= 8'hFF;
            13'd5154: data <= 8'h80;
            13'd5155: data <= 8'h00;
            13'd5156: data <= 8'h00;
            13'd5157: data <= 8'h00;
            13'd5158: data <= 8'h00;
            13'd5159: data <= 8'h00;
            13'd5160: data <= 8'h00;
            13'd5161: data <= 8'h00;
            13'd5162: data <= 8'h00;
            13'd5163: data <= 8'h00;
            13'd5164: data <= 8'h00;
            13'd5165: data <= 8'h03;
            13'd5166: data <= 8'hFF;
            13'd5167: data <= 8'hE1;
            13'd5168: data <= 8'hFE;
            13'd5169: data <= 8'h38;
            13'd5170: data <= 8'hFF;
            13'd5171: data <= 8'h8F;
            13'd5172: data <= 8'hFF;
            13'd5173: data <= 8'hFE;
            13'd5174: data <= 8'h00;
            13'd5175: data <= 8'h00;
            13'd5176: data <= 8'hFF;
            13'd5177: data <= 8'hFB;
            13'd5178: data <= 8'hFF;
            13'd5179: data <= 8'hFE;
            13'd5180: data <= 8'hFF;
            13'd5181: data <= 8'hFC;
            13'd5182: data <= 8'h1F;
            13'd5183: data <= 8'hFF;
            13'd5184: data <= 8'h80;
            13'd5185: data <= 8'h00;
            13'd5186: data <= 8'h00;
            13'd5187: data <= 8'h00;
            13'd5188: data <= 8'h00;
            13'd5189: data <= 8'h00;
            13'd5190: data <= 8'h00;
            13'd5191: data <= 8'h00;
            13'd5192: data <= 8'h00;
            13'd5193: data <= 8'h00;
            13'd5194: data <= 8'h00;
            13'd5195: data <= 8'h03;
            13'd5196: data <= 8'hFF;
            13'd5197: data <= 8'hFF;
            13'd5198: data <= 8'hFF;
            13'd5199: data <= 8'hFF;
            13'd5200: data <= 8'hFF;
            13'd5201: data <= 8'hFF;
            13'd5202: data <= 8'hFF;
            13'd5203: data <= 8'hFF;
            13'd5204: data <= 8'hFF;
            13'd5205: data <= 8'hFF;
            13'd5206: data <= 8'hFF;
            13'd5207: data <= 8'hBD;
            13'd5208: data <= 8'hFF;
            13'd5209: data <= 8'hFE;
            13'd5210: data <= 8'hFF;
            13'd5211: data <= 8'hFF;
            13'd5212: data <= 8'hFF;
            13'd5213: data <= 8'hFF;
            13'd5214: data <= 8'h80;
            13'd5215: data <= 8'h00;
            13'd5216: data <= 8'h00;
            13'd5217: data <= 8'h00;
            13'd5218: data <= 8'h00;
            13'd5219: data <= 8'h00;
            13'd5220: data <= 8'h00;
            13'd5221: data <= 8'h00;
            13'd5222: data <= 8'h00;
            13'd5223: data <= 8'h00;
            13'd5224: data <= 8'h00;
            13'd5225: data <= 8'h03;
            13'd5226: data <= 8'hFF;
            13'd5227: data <= 8'hFF;
            13'd5228: data <= 8'hFF;
            13'd5229: data <= 8'hFF;
            13'd5230: data <= 8'hFF;
            13'd5231: data <= 8'hFF;
            13'd5232: data <= 8'hFF;
            13'd5233: data <= 8'hFF;
            13'd5234: data <= 8'hFF;
            13'd5235: data <= 8'hFF;
            13'd5236: data <= 8'hFF;
            13'd5237: data <= 8'hBE;
            13'd5238: data <= 8'h7F;
            13'd5239: data <= 8'hFE;
            13'd5240: data <= 8'h7F;
            13'd5241: data <= 8'hFF;
            13'd5242: data <= 8'hFF;
            13'd5243: data <= 8'hFF;
            13'd5244: data <= 8'h80;
            13'd5245: data <= 8'h00;
            13'd5246: data <= 8'h00;
            13'd5247: data <= 8'h00;
            13'd5248: data <= 8'h00;
            13'd5249: data <= 8'h00;
            13'd5250: data <= 8'h00;
            13'd5251: data <= 8'h00;
            13'd5252: data <= 8'h00;
            13'd5253: data <= 8'h00;
            13'd5254: data <= 8'h00;
            13'd5255: data <= 8'h03;
            13'd5256: data <= 8'hFF;
            13'd5257: data <= 8'hFF;
            13'd5258: data <= 8'hFF;
            13'd5259: data <= 8'hFF;
            13'd5260: data <= 8'hFF;
            13'd5261: data <= 8'hFF;
            13'd5262: data <= 8'hFF;
            13'd5263: data <= 8'hFF;
            13'd5264: data <= 8'hFF;
            13'd5265: data <= 8'hFF;
            13'd5266: data <= 8'hFF;
            13'd5267: data <= 8'hBF;
            13'd5268: data <= 8'h03;
            13'd5269: data <= 8'hFE;
            13'd5270: data <= 8'h7F;
            13'd5271: data <= 8'hFF;
            13'd5272: data <= 8'hFF;
            13'd5273: data <= 8'hFF;
            13'd5274: data <= 8'h80;
            13'd5275: data <= 8'h00;
            13'd5276: data <= 8'h00;
            13'd5277: data <= 8'h00;
            13'd5278: data <= 8'h00;
            13'd5279: data <= 8'h00;
            13'd5280: data <= 8'h00;
            13'd5281: data <= 8'h00;
            13'd5282: data <= 8'h00;
            13'd5283: data <= 8'h00;
            13'd5284: data <= 8'h00;
            13'd5285: data <= 8'h03;
            13'd5286: data <= 8'hFF;
            13'd5287: data <= 8'hFF;
            13'd5288: data <= 8'hFF;
            13'd5289: data <= 8'hFF;
            13'd5290: data <= 8'hFF;
            13'd5291: data <= 8'hFF;
            13'd5292: data <= 8'hFF;
            13'd5293: data <= 8'hFF;
            13'd5294: data <= 8'hFF;
            13'd5295: data <= 8'hFF;
            13'd5296: data <= 8'hFF;
            13'd5297: data <= 8'hBF;
            13'd5298: data <= 8'hFF;
            13'd5299: data <= 8'hFF;
            13'd5300: data <= 8'h7F;
            13'd5301: data <= 8'hFF;
            13'd5302: data <= 8'hFF;
            13'd5303: data <= 8'hFF;
            13'd5304: data <= 8'h80;
            13'd5305: data <= 8'h00;
            13'd5306: data <= 8'h00;
            13'd5307: data <= 8'h00;
            13'd5308: data <= 8'h00;
            13'd5309: data <= 8'h00;
            13'd5310: data <= 8'h00;
            13'd5311: data <= 8'h00;
            13'd5312: data <= 8'h00;
            13'd5313: data <= 8'h00;
            13'd5314: data <= 8'h00;
            13'd5315: data <= 8'h03;
            13'd5316: data <= 8'hFF;
            13'd5317: data <= 8'hFF;
            13'd5318: data <= 8'hFF;
            13'd5319: data <= 8'hFF;
            13'd5320: data <= 8'hFF;
            13'd5321: data <= 8'hFF;
            13'd5322: data <= 8'hFF;
            13'd5323: data <= 8'hFF;
            13'd5324: data <= 8'hFF;
            13'd5325: data <= 8'hFF;
            13'd5326: data <= 8'hFF;
            13'd5327: data <= 8'hBF;
            13'd5328: data <= 8'hFF;
            13'd5329: data <= 8'hFF;
            13'd5330: data <= 8'h7F;
            13'd5331: data <= 8'hFF;
            13'd5332: data <= 8'hFF;
            13'd5333: data <= 8'hFF;
            13'd5334: data <= 8'h80;
            13'd5335: data <= 8'h00;
            13'd5336: data <= 8'h00;
            13'd5337: data <= 8'h00;
            13'd5338: data <= 8'h00;
            13'd5339: data <= 8'h00;
            13'd5340: data <= 8'h00;
            13'd5341: data <= 8'h00;
            13'd5342: data <= 8'h00;
            13'd5343: data <= 8'h00;
            13'd5344: data <= 8'h00;
            13'd5345: data <= 8'h03;
            13'd5346: data <= 8'hFF;
            13'd5347: data <= 8'hFF;
            13'd5348: data <= 8'hFF;
            13'd5349: data <= 8'hFF;
            13'd5350: data <= 8'hFF;
            13'd5351: data <= 8'hFF;
            13'd5352: data <= 8'hFF;
            13'd5353: data <= 8'hFF;
            13'd5354: data <= 8'hFF;
            13'd5355: data <= 8'hFF;
            13'd5356: data <= 8'hFF;
            13'd5357: data <= 8'hBF;
            13'd5358: data <= 8'hFF;
            13'd5359: data <= 8'hFF;
            13'd5360: data <= 8'hFF;
            13'd5361: data <= 8'hFF;
            13'd5362: data <= 8'hFF;
            13'd5363: data <= 8'hFF;
            13'd5364: data <= 8'h80;
            13'd5365: data <= 8'h00;
            13'd5366: data <= 8'h00;
            13'd5367: data <= 8'h00;
            13'd5368: data <= 8'h00;
            13'd5369: data <= 8'h00;
            13'd5370: data <= 8'h00;
            13'd5371: data <= 8'h00;
            13'd5372: data <= 8'h00;
            13'd5373: data <= 8'h00;
            13'd5374: data <= 8'h00;
            13'd5375: data <= 8'h03;
            13'd5376: data <= 8'hFF;
            13'd5377: data <= 8'hFF;
            13'd5378: data <= 8'hFF;
            13'd5379: data <= 8'hFF;
            13'd5380: data <= 8'hFF;
            13'd5381: data <= 8'hFF;
            13'd5382: data <= 8'hFF;
            13'd5383: data <= 8'hFF;
            13'd5384: data <= 8'hFF;
            13'd5385: data <= 8'hFF;
            13'd5386: data <= 8'hFF;
            13'd5387: data <= 8'hFF;
            13'd5388: data <= 8'hFF;
            13'd5389: data <= 8'hFF;
            13'd5390: data <= 8'hFF;
            13'd5391: data <= 8'hFF;
            13'd5392: data <= 8'hFF;
            13'd5393: data <= 8'hFF;
            13'd5394: data <= 8'h80;
            13'd5395: data <= 8'h00;
            13'd5396: data <= 8'h00;
            13'd5397: data <= 8'h00;
            13'd5398: data <= 8'h00;
            13'd5399: data <= 8'h00;
            default: data <= 8'h00;
        endcase
    end

endmodule
