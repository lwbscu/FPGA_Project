// ============================================================================
// Module: pic_ram
// Description: 图片RAM模块 - 存储简单的白色背景和球的图像数据
// Author: GitHub Copilot
// Date: 2025-05-28
// ============================================================================

`timescale 1 ns / 100 ps

module pic_ram (
    input wire [8:0] address,
    output reg [239:0] q,
    input wire [8:0] offset
);
      // 创建简单的白色背景和球的图案
    always @ (*) begin
        case(address - offset)
            // 球的图案（黑色球，使用0表示黑色像素，1表示白色背景）
            9'd1:   q = 240'h000000000000000000000FFFF800000000000000000000000000000000; // 球的顶部
            9'd2:   q = 240'h0000000000000000000FFFFFFF0000000000000000000000000000000; 
            9'd3:   q = 240'h000000000000000000FFFFFFFFF800000000000000000000000000000;
            9'd4:   q = 240'h000000000000000000FFFFFFFFF800000000000000000000000000000;
            9'd5:   q = 240'h00000000000000000FFFFFFFFFFF00000000000000000000000000000; // 球的中部（最宽）
            9'd6:   q = 240'h00000000000000000FFFFFFFFFFF00000000000000000000000000000;
            9'd7:   q = 240'h000000000000000000FFFFFFFFF800000000000000000000000000000;
            9'd8:   q = 240'h000000000000000000FFFFFFFFF800000000000000000000000000000;
            9'd9:   q = 240'h0000000000000000000FFFFFFF0000000000000000000000000000000;
            9'd10:  q = 240'h000000000000000000000FFFF800000000000000000000000000000000; // 球的底部
            
            // 添加手柄线条（水平线，黑色）
            9'd200: q = 240'h000000000000000000000000000000000000000000000000000000000000; // 全黑水平线
            9'd201: q = 240'h000000000000000000000000000000000000000000000000000000000000; // 全黑水平线
            9'd202: q = 240'h000000000000000000000000000000000000000000000000000000000000; // 全黑水平线
            
            // 为了测试显示，添加更多可见图案
            9'd50:  q = 240'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA; // 棋盘格图案
            9'd51:  q = 240'h555555555555555555555555555555555555555555555555555555555555; // 反相棋盘格
            9'd52:  q = 240'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA; // 棋盘格图案
            
            // 边界线条测试
            9'd100: q = 240'h000000000000000000000000000000000000000000000000000000000000; // 全黑线
            9'd300: q = 240'h000000000000000000000000000000000000000000000000000000000000; // 全黑线
            
            // 默认为白色背景（1表示白色像素）
            default: q = 240'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF; // 白色背景
        endcase
    end

endmodule
