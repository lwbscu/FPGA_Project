// �Զ����ɵ�ROMģ��
// ͼƬ�ߴ�: 120 x 160
// ��ɫ��ʽ: RGB565(16λ)
// ���ݴ�С: 38400 �ֽ�

module test_pattern_rom (
    input wire clk,
    input wire [15:0] addr,
    output reg [7:0] data
);

    // ROM���ݴ洢 (38400 ����ַ)
    always @(posedge clk) begin
        case (addr)
            16'd0: data <= 8'hFF;
            16'd1: data <= 8'hFF;
            16'd2: data <= 8'hFF;
            16'd3: data <= 8'hFF;
            16'd4: data <= 8'hFF;
            16'd5: data <= 8'hFF;
            16'd6: data <= 8'hFF;
            16'd7: data <= 8'hFF;
            16'd8: data <= 8'hFF;
            16'd9: data <= 8'hFF;
            16'd10: data <= 8'hFF;
            16'd11: data <= 8'hFF;
            16'd12: data <= 8'hFF;
            16'd13: data <= 8'hFF;
            16'd14: data <= 8'hFF;
            16'd15: data <= 8'hFF;
            16'd16: data <= 8'hFF;
            16'd17: data <= 8'hFF;
            16'd18: data <= 8'hFF;
            16'd19: data <= 8'hFF;
            16'd20: data <= 8'hFF;
            16'd21: data <= 8'hFF;
            16'd22: data <= 8'hFF;
            16'd23: data <= 8'hFF;
            16'd24: data <= 8'hFF;
            16'd25: data <= 8'hFF;
            16'd26: data <= 8'hFF;
            16'd27: data <= 8'hFF;
            16'd28: data <= 8'hFF;
            16'd29: data <= 8'hFF;
            16'd30: data <= 8'hFF;
            16'd31: data <= 8'hFF;
            16'd32: data <= 8'hFF;
            16'd33: data <= 8'hFF;
            16'd34: data <= 8'hFF;
            16'd35: data <= 8'hFF;
            16'd36: data <= 8'hFF;
            16'd37: data <= 8'hFF;
            16'd38: data <= 8'hFF;
            16'd39: data <= 8'hFF;
            16'd40: data <= 8'hFF;
            16'd41: data <= 8'hFF;
            16'd42: data <= 8'hFF;
            16'd43: data <= 8'hFF;
            16'd44: data <= 8'hFF;
            16'd45: data <= 8'hFF;
            16'd46: data <= 8'hFF;
            16'd47: data <= 8'hFF;
            16'd48: data <= 8'hFF;
            16'd49: data <= 8'hFF;
            16'd50: data <= 8'hFF;
            16'd51: data <= 8'hFF;
            16'd52: data <= 8'hFF;
            16'd53: data <= 8'hFF;
            16'd54: data <= 8'hFF;
            16'd55: data <= 8'hFF;
            16'd56: data <= 8'hFF;
            16'd57: data <= 8'hFF;
            16'd58: data <= 8'hFF;
            16'd59: data <= 8'hFF;
            16'd60: data <= 8'hFF;
            16'd61: data <= 8'hFF;
            16'd62: data <= 8'hFF;
            16'd63: data <= 8'hFF;
            16'd64: data <= 8'hFF;
            16'd65: data <= 8'hFF;
            16'd66: data <= 8'hFF;
            16'd67: data <= 8'hFF;
            16'd68: data <= 8'hFF;
            16'd69: data <= 8'hFF;
            16'd70: data <= 8'hFF;
            16'd71: data <= 8'hFF;
            16'd72: data <= 8'hFF;
            16'd73: data <= 8'hFF;
            16'd74: data <= 8'hFF;
            16'd75: data <= 8'hFF;
            16'd76: data <= 8'hFF;
            16'd77: data <= 8'hFF;
            16'd78: data <= 8'hFF;
            16'd79: data <= 8'hFF;
            16'd80: data <= 8'hFF;
            16'd81: data <= 8'hFF;
            16'd82: data <= 8'hFF;
            16'd83: data <= 8'hFF;
            16'd84: data <= 8'hFF;
            16'd85: data <= 8'hFF;
            16'd86: data <= 8'hFF;
            16'd87: data <= 8'hFF;
            16'd88: data <= 8'hFF;
            16'd89: data <= 8'hFF;
            16'd90: data <= 8'hFF;
            16'd91: data <= 8'hFF;
            16'd92: data <= 8'hFF;
            16'd93: data <= 8'hFF;
            16'd94: data <= 8'hFF;
            16'd95: data <= 8'hFF;
            16'd96: data <= 8'hFF;
            16'd97: data <= 8'hFF;
            16'd98: data <= 8'hFF;
            16'd99: data <= 8'hFF;
            16'd100: data <= 8'hFF;
            16'd101: data <= 8'hFF;
            16'd102: data <= 8'hFF;
            16'd103: data <= 8'hFF;
            16'd104: data <= 8'hFF;
            16'd105: data <= 8'hFF;
            16'd106: data <= 8'hFF;
            16'd107: data <= 8'hFF;
            16'd108: data <= 8'hFF;
            16'd109: data <= 8'hFF;
            16'd110: data <= 8'hFF;
            16'd111: data <= 8'hFF;
            16'd112: data <= 8'hFF;
            16'd113: data <= 8'hFF;
            16'd114: data <= 8'hFF;
            16'd115: data <= 8'hFF;
            16'd116: data <= 8'hFF;
            16'd117: data <= 8'hFF;
            16'd118: data <= 8'hFF;
            16'd119: data <= 8'hFF;
            16'd120: data <= 8'hFF;
            16'd121: data <= 8'hFF;
            16'd122: data <= 8'hFF;
            16'd123: data <= 8'hFF;
            16'd124: data <= 8'hFF;
            16'd125: data <= 8'hFF;
            16'd126: data <= 8'hFF;
            16'd127: data <= 8'hFF;
            16'd128: data <= 8'hFF;
            16'd129: data <= 8'hFF;
            16'd130: data <= 8'hFF;
            16'd131: data <= 8'hFF;
            16'd132: data <= 8'hFF;
            16'd133: data <= 8'hFF;
            16'd134: data <= 8'hFF;
            16'd135: data <= 8'hFF;
            16'd136: data <= 8'hFF;
            16'd137: data <= 8'hFF;
            16'd138: data <= 8'hFF;
            16'd139: data <= 8'hFF;
            16'd140: data <= 8'hFF;
            16'd141: data <= 8'hFF;
            16'd142: data <= 8'hFF;
            16'd143: data <= 8'hFF;
            16'd144: data <= 8'hFF;
            16'd145: data <= 8'hFF;
            16'd146: data <= 8'hFF;
            16'd147: data <= 8'hFF;
            16'd148: data <= 8'hFF;
            16'd149: data <= 8'hFF;
            16'd150: data <= 8'hFF;
            16'd151: data <= 8'hFF;
            16'd152: data <= 8'hFF;
            16'd153: data <= 8'hFF;
            16'd154: data <= 8'hFF;
            16'd155: data <= 8'hFF;
            16'd156: data <= 8'hFF;
            16'd157: data <= 8'hFF;
            16'd158: data <= 8'hFF;
            16'd159: data <= 8'hFF;
            16'd160: data <= 8'hFF;
            16'd161: data <= 8'hFF;
            16'd162: data <= 8'hFF;
            16'd163: data <= 8'hFF;
            16'd164: data <= 8'hFF;
            16'd165: data <= 8'hFF;
            16'd166: data <= 8'hFF;
            16'd167: data <= 8'hFF;
            16'd168: data <= 8'hFF;
            16'd169: data <= 8'hFF;
            16'd170: data <= 8'hFF;
            16'd171: data <= 8'hFF;
            16'd172: data <= 8'hFF;
            16'd173: data <= 8'hFF;
            16'd174: data <= 8'hFF;
            16'd175: data <= 8'hFF;
            16'd176: data <= 8'hFF;
            16'd177: data <= 8'hFF;
            16'd178: data <= 8'hFF;
            16'd179: data <= 8'hFF;
            16'd180: data <= 8'hFF;
            16'd181: data <= 8'hFF;
            16'd182: data <= 8'hFF;
            16'd183: data <= 8'hFF;
            16'd184: data <= 8'hFF;
            16'd185: data <= 8'hFF;
            16'd186: data <= 8'hFF;
            16'd187: data <= 8'hFF;
            16'd188: data <= 8'hFF;
            16'd189: data <= 8'hFF;
            16'd190: data <= 8'hFF;
            16'd191: data <= 8'hFF;
            16'd192: data <= 8'hFF;
            16'd193: data <= 8'hFF;
            16'd194: data <= 8'hFF;
            16'd195: data <= 8'hFF;
            16'd196: data <= 8'hFF;
            16'd197: data <= 8'hFF;
            16'd198: data <= 8'hFF;
            16'd199: data <= 8'hFF;
            16'd200: data <= 8'hFF;
            16'd201: data <= 8'hFF;
            16'd202: data <= 8'hFF;
            16'd203: data <= 8'hFF;
            16'd204: data <= 8'hFF;
            16'd205: data <= 8'hFF;
            16'd206: data <= 8'hFF;
            16'd207: data <= 8'hFF;
            16'd208: data <= 8'hFF;
            16'd209: data <= 8'hFF;
            16'd210: data <= 8'hFF;
            16'd211: data <= 8'hFF;
            16'd212: data <= 8'hFF;
            16'd213: data <= 8'hFF;
            16'd214: data <= 8'hFF;
            16'd215: data <= 8'hFF;
            16'd216: data <= 8'hFF;
            16'd217: data <= 8'hFF;
            16'd218: data <= 8'hFF;
            16'd219: data <= 8'hFF;
            16'd220: data <= 8'hFF;
            16'd221: data <= 8'hFF;
            16'd222: data <= 8'hFF;
            16'd223: data <= 8'hFF;
            16'd224: data <= 8'hFF;
            16'd225: data <= 8'hFF;
            16'd226: data <= 8'hFF;
            16'd227: data <= 8'hFF;
            16'd228: data <= 8'hFF;
            16'd229: data <= 8'hFF;
            16'd230: data <= 8'hFF;
            16'd231: data <= 8'hFF;
            16'd232: data <= 8'hFF;
            16'd233: data <= 8'hFF;
            16'd234: data <= 8'hFF;
            16'd235: data <= 8'hFF;
            16'd236: data <= 8'hFF;
            16'd237: data <= 8'hFF;
            16'd238: data <= 8'hFF;
            16'd239: data <= 8'hFF;
            16'd240: data <= 8'hFF;
            16'd241: data <= 8'hFF;
            16'd242: data <= 8'h00;
            16'd243: data <= 8'hF8;
            16'd244: data <= 8'h00;
            16'd245: data <= 8'hF8;
            16'd246: data <= 8'h00;
            16'd247: data <= 8'hF8;
            16'd248: data <= 8'h00;
            16'd249: data <= 8'hF8;
            16'd250: data <= 8'h00;
            16'd251: data <= 8'hF8;
            16'd252: data <= 8'h00;
            16'd253: data <= 8'hF8;
            16'd254: data <= 8'h00;
            16'd255: data <= 8'hF8;
            16'd256: data <= 8'h00;
            16'd257: data <= 8'hF8;
            16'd258: data <= 8'h00;
            16'd259: data <= 8'hF8;
            16'd260: data <= 8'h00;
            16'd261: data <= 8'hF8;
            16'd262: data <= 8'h00;
            16'd263: data <= 8'hF8;
            16'd264: data <= 8'h00;
            16'd265: data <= 8'hF8;
            16'd266: data <= 8'h00;
            16'd267: data <= 8'hF8;
            16'd268: data <= 8'h00;
            16'd269: data <= 8'hF8;
            16'd270: data <= 8'h00;
            16'd271: data <= 8'hF8;
            16'd272: data <= 8'h00;
            16'd273: data <= 8'hF8;
            16'd274: data <= 8'h00;
            16'd275: data <= 8'hF8;
            16'd276: data <= 8'h00;
            16'd277: data <= 8'hF8;
            16'd278: data <= 8'h00;
            16'd279: data <= 8'hF8;
            16'd280: data <= 8'hFF;
            16'd281: data <= 8'hFF;
            16'd282: data <= 8'h00;
            16'd283: data <= 8'hF8;
            16'd284: data <= 8'h00;
            16'd285: data <= 8'hF8;
            16'd286: data <= 8'h00;
            16'd287: data <= 8'hF8;
            16'd288: data <= 8'h00;
            16'd289: data <= 8'hF8;
            16'd290: data <= 8'h00;
            16'd291: data <= 8'hF8;
            16'd292: data <= 8'h00;
            16'd293: data <= 8'hF8;
            16'd294: data <= 8'h00;
            16'd295: data <= 8'hF8;
            16'd296: data <= 8'h00;
            16'd297: data <= 8'hF8;
            16'd298: data <= 8'h00;
            16'd299: data <= 8'hF8;
            16'd300: data <= 8'h00;
            16'd301: data <= 8'hF8;
            16'd302: data <= 8'h00;
            16'd303: data <= 8'hF8;
            16'd304: data <= 8'h00;
            16'd305: data <= 8'hF8;
            16'd306: data <= 8'h00;
            16'd307: data <= 8'hF8;
            16'd308: data <= 8'h00;
            16'd309: data <= 8'hF8;
            16'd310: data <= 8'h00;
            16'd311: data <= 8'hF8;
            16'd312: data <= 8'h00;
            16'd313: data <= 8'hF8;
            16'd314: data <= 8'h00;
            16'd315: data <= 8'hF8;
            16'd316: data <= 8'h00;
            16'd317: data <= 8'hF8;
            16'd318: data <= 8'h00;
            16'd319: data <= 8'hF8;
            16'd320: data <= 8'hFF;
            16'd321: data <= 8'hFF;
            16'd322: data <= 8'h00;
            16'd323: data <= 8'hF8;
            16'd324: data <= 8'h00;
            16'd325: data <= 8'hF8;
            16'd326: data <= 8'h00;
            16'd327: data <= 8'hF8;
            16'd328: data <= 8'h00;
            16'd329: data <= 8'hF8;
            16'd330: data <= 8'h00;
            16'd331: data <= 8'hF8;
            16'd332: data <= 8'h00;
            16'd333: data <= 8'hF8;
            16'd334: data <= 8'h00;
            16'd335: data <= 8'hF8;
            16'd336: data <= 8'h00;
            16'd337: data <= 8'hF8;
            16'd338: data <= 8'h00;
            16'd339: data <= 8'hF8;
            16'd340: data <= 8'h00;
            16'd341: data <= 8'hF8;
            16'd342: data <= 8'h00;
            16'd343: data <= 8'hF8;
            16'd344: data <= 8'h00;
            16'd345: data <= 8'hF8;
            16'd346: data <= 8'h00;
            16'd347: data <= 8'hF8;
            16'd348: data <= 8'h00;
            16'd349: data <= 8'hF8;
            16'd350: data <= 8'h00;
            16'd351: data <= 8'hF8;
            16'd352: data <= 8'h00;
            16'd353: data <= 8'hF8;
            16'd354: data <= 8'h00;
            16'd355: data <= 8'hF8;
            16'd356: data <= 8'h00;
            16'd357: data <= 8'hF8;
            16'd358: data <= 8'h00;
            16'd359: data <= 8'hF8;
            16'd360: data <= 8'hFF;
            16'd361: data <= 8'hFF;
            16'd362: data <= 8'h00;
            16'd363: data <= 8'hF8;
            16'd364: data <= 8'h00;
            16'd365: data <= 8'hF8;
            16'd366: data <= 8'h00;
            16'd367: data <= 8'hF8;
            16'd368: data <= 8'h00;
            16'd369: data <= 8'hF8;
            16'd370: data <= 8'h00;
            16'd371: data <= 8'hF8;
            16'd372: data <= 8'h00;
            16'd373: data <= 8'hF8;
            16'd374: data <= 8'h00;
            16'd375: data <= 8'hF8;
            16'd376: data <= 8'h00;
            16'd377: data <= 8'hF8;
            16'd378: data <= 8'h00;
            16'd379: data <= 8'hF8;
            16'd380: data <= 8'h00;
            16'd381: data <= 8'hF8;
            16'd382: data <= 8'h00;
            16'd383: data <= 8'hF8;
            16'd384: data <= 8'h00;
            16'd385: data <= 8'hF8;
            16'd386: data <= 8'h00;
            16'd387: data <= 8'hF8;
            16'd388: data <= 8'h00;
            16'd389: data <= 8'hF8;
            16'd390: data <= 8'h00;
            16'd391: data <= 8'hF8;
            16'd392: data <= 8'h00;
            16'd393: data <= 8'hF8;
            16'd394: data <= 8'h00;
            16'd395: data <= 8'hF8;
            16'd396: data <= 8'h00;
            16'd397: data <= 8'hF8;
            16'd398: data <= 8'h00;
            16'd399: data <= 8'hF8;
            16'd400: data <= 8'hFF;
            16'd401: data <= 8'hFF;
            16'd402: data <= 8'h00;
            16'd403: data <= 8'hF8;
            16'd404: data <= 8'h00;
            16'd405: data <= 8'hF8;
            16'd406: data <= 8'h00;
            16'd407: data <= 8'hF8;
            16'd408: data <= 8'h00;
            16'd409: data <= 8'hF8;
            16'd410: data <= 8'h00;
            16'd411: data <= 8'hF8;
            16'd412: data <= 8'h00;
            16'd413: data <= 8'hF8;
            16'd414: data <= 8'h00;
            16'd415: data <= 8'hF8;
            16'd416: data <= 8'h00;
            16'd417: data <= 8'hF8;
            16'd418: data <= 8'h00;
            16'd419: data <= 8'hF8;
            16'd420: data <= 8'h00;
            16'd421: data <= 8'hF8;
            16'd422: data <= 8'h00;
            16'd423: data <= 8'hF8;
            16'd424: data <= 8'h00;
            16'd425: data <= 8'hF8;
            16'd426: data <= 8'h00;
            16'd427: data <= 8'hF8;
            16'd428: data <= 8'h00;
            16'd429: data <= 8'hF8;
            16'd430: data <= 8'h00;
            16'd431: data <= 8'hF8;
            16'd432: data <= 8'h00;
            16'd433: data <= 8'hF8;
            16'd434: data <= 8'h00;
            16'd435: data <= 8'hF8;
            16'd436: data <= 8'h00;
            16'd437: data <= 8'hF8;
            16'd438: data <= 8'h00;
            16'd439: data <= 8'hF8;
            16'd440: data <= 8'hFF;
            16'd441: data <= 8'hFF;
            16'd442: data <= 8'h00;
            16'd443: data <= 8'hF8;
            16'd444: data <= 8'h00;
            16'd445: data <= 8'hF8;
            16'd446: data <= 8'h00;
            16'd447: data <= 8'hF8;
            16'd448: data <= 8'h00;
            16'd449: data <= 8'hF8;
            16'd450: data <= 8'h00;
            16'd451: data <= 8'hF8;
            16'd452: data <= 8'h00;
            16'd453: data <= 8'hF8;
            16'd454: data <= 8'h00;
            16'd455: data <= 8'hF8;
            16'd456: data <= 8'h00;
            16'd457: data <= 8'hF8;
            16'd458: data <= 8'h00;
            16'd459: data <= 8'hF8;
            16'd460: data <= 8'h00;
            16'd461: data <= 8'hF8;
            16'd462: data <= 8'h00;
            16'd463: data <= 8'hF8;
            16'd464: data <= 8'h00;
            16'd465: data <= 8'hF8;
            16'd466: data <= 8'h00;
            16'd467: data <= 8'hF8;
            16'd468: data <= 8'h00;
            16'd469: data <= 8'hF8;
            16'd470: data <= 8'h00;
            16'd471: data <= 8'hF8;
            16'd472: data <= 8'h00;
            16'd473: data <= 8'hF8;
            16'd474: data <= 8'h00;
            16'd475: data <= 8'hF8;
            16'd476: data <= 8'h00;
            16'd477: data <= 8'hF8;
            16'd478: data <= 8'h00;
            16'd479: data <= 8'hF8;
            16'd480: data <= 8'hFF;
            16'd481: data <= 8'hFF;
            16'd482: data <= 8'h00;
            16'd483: data <= 8'hF8;
            16'd484: data <= 8'h00;
            16'd485: data <= 8'hF8;
            16'd486: data <= 8'h00;
            16'd487: data <= 8'hF8;
            16'd488: data <= 8'h00;
            16'd489: data <= 8'hF8;
            16'd490: data <= 8'h00;
            16'd491: data <= 8'hF8;
            16'd492: data <= 8'h00;
            16'd493: data <= 8'hF8;
            16'd494: data <= 8'h00;
            16'd495: data <= 8'hF8;
            16'd496: data <= 8'h00;
            16'd497: data <= 8'hF8;
            16'd498: data <= 8'h00;
            16'd499: data <= 8'hF8;
            16'd500: data <= 8'h00;
            16'd501: data <= 8'hF8;
            16'd502: data <= 8'h00;
            16'd503: data <= 8'hF8;
            16'd504: data <= 8'h00;
            16'd505: data <= 8'hF8;
            16'd506: data <= 8'h00;
            16'd507: data <= 8'hF8;
            16'd508: data <= 8'h00;
            16'd509: data <= 8'hF8;
            16'd510: data <= 8'h00;
            16'd511: data <= 8'hF8;
            16'd512: data <= 8'h00;
            16'd513: data <= 8'hF8;
            16'd514: data <= 8'h00;
            16'd515: data <= 8'hF8;
            16'd516: data <= 8'h00;
            16'd517: data <= 8'hF8;
            16'd518: data <= 8'h00;
            16'd519: data <= 8'hF8;
            16'd520: data <= 8'hFF;
            16'd521: data <= 8'hFF;
            16'd522: data <= 8'h00;
            16'd523: data <= 8'hF8;
            16'd524: data <= 8'h00;
            16'd525: data <= 8'hF8;
            16'd526: data <= 8'h00;
            16'd527: data <= 8'hF8;
            16'd528: data <= 8'h00;
            16'd529: data <= 8'hF8;
            16'd530: data <= 8'h00;
            16'd531: data <= 8'hF8;
            16'd532: data <= 8'h00;
            16'd533: data <= 8'hF8;
            16'd534: data <= 8'h00;
            16'd535: data <= 8'hF8;
            16'd536: data <= 8'h00;
            16'd537: data <= 8'hF8;
            16'd538: data <= 8'h00;
            16'd539: data <= 8'hF8;
            16'd540: data <= 8'h00;
            16'd541: data <= 8'hF8;
            16'd542: data <= 8'h00;
            16'd543: data <= 8'hF8;
            16'd544: data <= 8'h00;
            16'd545: data <= 8'hF8;
            16'd546: data <= 8'h00;
            16'd547: data <= 8'hF8;
            16'd548: data <= 8'h00;
            16'd549: data <= 8'hF8;
            16'd550: data <= 8'h00;
            16'd551: data <= 8'hF8;
            16'd552: data <= 8'h00;
            16'd553: data <= 8'hF8;
            16'd554: data <= 8'h00;
            16'd555: data <= 8'hF8;
            16'd556: data <= 8'h00;
            16'd557: data <= 8'hF8;
            16'd558: data <= 8'h00;
            16'd559: data <= 8'hF8;
            16'd560: data <= 8'hFF;
            16'd561: data <= 8'hFF;
            16'd562: data <= 8'h00;
            16'd563: data <= 8'hF8;
            16'd564: data <= 8'h00;
            16'd565: data <= 8'hF8;
            16'd566: data <= 8'h00;
            16'd567: data <= 8'hF8;
            16'd568: data <= 8'h00;
            16'd569: data <= 8'hF8;
            16'd570: data <= 8'h00;
            16'd571: data <= 8'hF8;
            16'd572: data <= 8'h00;
            16'd573: data <= 8'hF8;
            16'd574: data <= 8'h00;
            16'd575: data <= 8'hF8;
            16'd576: data <= 8'h00;
            16'd577: data <= 8'hF8;
            16'd578: data <= 8'h00;
            16'd579: data <= 8'hF8;
            16'd580: data <= 8'h00;
            16'd581: data <= 8'hF8;
            16'd582: data <= 8'h00;
            16'd583: data <= 8'hF8;
            16'd584: data <= 8'h00;
            16'd585: data <= 8'hF8;
            16'd586: data <= 8'h00;
            16'd587: data <= 8'hF8;
            16'd588: data <= 8'h00;
            16'd589: data <= 8'hF8;
            16'd590: data <= 8'h00;
            16'd591: data <= 8'hF8;
            16'd592: data <= 8'h00;
            16'd593: data <= 8'hF8;
            16'd594: data <= 8'h00;
            16'd595: data <= 8'hF8;
            16'd596: data <= 8'h00;
            16'd597: data <= 8'hF8;
            16'd598: data <= 8'h00;
            16'd599: data <= 8'hF8;
            16'd600: data <= 8'hFF;
            16'd601: data <= 8'hFF;
            16'd602: data <= 8'h00;
            16'd603: data <= 8'hF8;
            16'd604: data <= 8'h00;
            16'd605: data <= 8'hF8;
            16'd606: data <= 8'h00;
            16'd607: data <= 8'hF8;
            16'd608: data <= 8'h00;
            16'd609: data <= 8'hF8;
            16'd610: data <= 8'h00;
            16'd611: data <= 8'hF8;
            16'd612: data <= 8'h00;
            16'd613: data <= 8'hF8;
            16'd614: data <= 8'h00;
            16'd615: data <= 8'hF8;
            16'd616: data <= 8'h00;
            16'd617: data <= 8'hF8;
            16'd618: data <= 8'h00;
            16'd619: data <= 8'hF8;
            16'd620: data <= 8'h00;
            16'd621: data <= 8'hF8;
            16'd622: data <= 8'h00;
            16'd623: data <= 8'hF8;
            16'd624: data <= 8'h00;
            16'd625: data <= 8'hF8;
            16'd626: data <= 8'h00;
            16'd627: data <= 8'hF8;
            16'd628: data <= 8'h00;
            16'd629: data <= 8'hF8;
            16'd630: data <= 8'h00;
            16'd631: data <= 8'hF8;
            16'd632: data <= 8'h00;
            16'd633: data <= 8'hF8;
            16'd634: data <= 8'h00;
            16'd635: data <= 8'hF8;
            16'd636: data <= 8'h00;
            16'd637: data <= 8'hF8;
            16'd638: data <= 8'h00;
            16'd639: data <= 8'hF8;
            16'd640: data <= 8'hFF;
            16'd641: data <= 8'hFF;
            16'd642: data <= 8'h00;
            16'd643: data <= 8'hF8;
            16'd644: data <= 8'h00;
            16'd645: data <= 8'hF8;
            16'd646: data <= 8'h00;
            16'd647: data <= 8'hF8;
            16'd648: data <= 8'h00;
            16'd649: data <= 8'hF8;
            16'd650: data <= 8'h00;
            16'd651: data <= 8'hF8;
            16'd652: data <= 8'h00;
            16'd653: data <= 8'hF8;
            16'd654: data <= 8'h00;
            16'd655: data <= 8'hF8;
            16'd656: data <= 8'h00;
            16'd657: data <= 8'hF8;
            16'd658: data <= 8'h00;
            16'd659: data <= 8'hF8;
            16'd660: data <= 8'h00;
            16'd661: data <= 8'hF8;
            16'd662: data <= 8'h00;
            16'd663: data <= 8'hF8;
            16'd664: data <= 8'h00;
            16'd665: data <= 8'hF8;
            16'd666: data <= 8'h00;
            16'd667: data <= 8'hF8;
            16'd668: data <= 8'h00;
            16'd669: data <= 8'hF8;
            16'd670: data <= 8'h00;
            16'd671: data <= 8'hF8;
            16'd672: data <= 8'h00;
            16'd673: data <= 8'hF8;
            16'd674: data <= 8'h00;
            16'd675: data <= 8'hF8;
            16'd676: data <= 8'h00;
            16'd677: data <= 8'hF8;
            16'd678: data <= 8'h00;
            16'd679: data <= 8'hF8;
            16'd680: data <= 8'hFF;
            16'd681: data <= 8'hFF;
            16'd682: data <= 8'h00;
            16'd683: data <= 8'hF8;
            16'd684: data <= 8'h00;
            16'd685: data <= 8'hF8;
            16'd686: data <= 8'h00;
            16'd687: data <= 8'hF8;
            16'd688: data <= 8'h00;
            16'd689: data <= 8'hF8;
            16'd690: data <= 8'h00;
            16'd691: data <= 8'hF8;
            16'd692: data <= 8'h00;
            16'd693: data <= 8'hF8;
            16'd694: data <= 8'h00;
            16'd695: data <= 8'hF8;
            16'd696: data <= 8'h00;
            16'd697: data <= 8'hF8;
            16'd698: data <= 8'h00;
            16'd699: data <= 8'hF8;
            16'd700: data <= 8'h00;
            16'd701: data <= 8'hF8;
            16'd702: data <= 8'h00;
            16'd703: data <= 8'hF8;
            16'd704: data <= 8'h00;
            16'd705: data <= 8'hF8;
            16'd706: data <= 8'h00;
            16'd707: data <= 8'hF8;
            16'd708: data <= 8'h00;
            16'd709: data <= 8'hF8;
            16'd710: data <= 8'h00;
            16'd711: data <= 8'hF8;
            16'd712: data <= 8'h00;
            16'd713: data <= 8'hF8;
            16'd714: data <= 8'h00;
            16'd715: data <= 8'hF8;
            16'd716: data <= 8'h00;
            16'd717: data <= 8'hF8;
            16'd718: data <= 8'h00;
            16'd719: data <= 8'hF8;
            16'd720: data <= 8'hFF;
            16'd721: data <= 8'hFF;
            16'd722: data <= 8'h00;
            16'd723: data <= 8'hF8;
            16'd724: data <= 8'h00;
            16'd725: data <= 8'hF8;
            16'd726: data <= 8'h00;
            16'd727: data <= 8'hF8;
            16'd728: data <= 8'h00;
            16'd729: data <= 8'hF8;
            16'd730: data <= 8'h00;
            16'd731: data <= 8'hF8;
            16'd732: data <= 8'h00;
            16'd733: data <= 8'hF8;
            16'd734: data <= 8'h00;
            16'd735: data <= 8'hF8;
            16'd736: data <= 8'h00;
            16'd737: data <= 8'hF8;
            16'd738: data <= 8'h00;
            16'd739: data <= 8'hF8;
            16'd740: data <= 8'h00;
            16'd741: data <= 8'hF8;
            16'd742: data <= 8'h00;
            16'd743: data <= 8'hF8;
            16'd744: data <= 8'h00;
            16'd745: data <= 8'hF8;
            16'd746: data <= 8'h00;
            16'd747: data <= 8'hF8;
            16'd748: data <= 8'h00;
            16'd749: data <= 8'hF8;
            16'd750: data <= 8'h00;
            16'd751: data <= 8'hF8;
            16'd752: data <= 8'h00;
            16'd753: data <= 8'hF8;
            16'd754: data <= 8'h00;
            16'd755: data <= 8'hF8;
            16'd756: data <= 8'h00;
            16'd757: data <= 8'hF8;
            16'd758: data <= 8'h00;
            16'd759: data <= 8'hF8;
            16'd760: data <= 8'hFF;
            16'd761: data <= 8'hFF;
            16'd762: data <= 8'h00;
            16'd763: data <= 8'hF8;
            16'd764: data <= 8'h00;
            16'd765: data <= 8'hF8;
            16'd766: data <= 8'h00;
            16'd767: data <= 8'hF8;
            16'd768: data <= 8'h00;
            16'd769: data <= 8'hF8;
            16'd770: data <= 8'h00;
            16'd771: data <= 8'hF8;
            16'd772: data <= 8'h00;
            16'd773: data <= 8'hF8;
            16'd774: data <= 8'h00;
            16'd775: data <= 8'hF8;
            16'd776: data <= 8'h00;
            16'd777: data <= 8'hF8;
            16'd778: data <= 8'h00;
            16'd779: data <= 8'hF8;
            16'd780: data <= 8'h00;
            16'd781: data <= 8'hF8;
            16'd782: data <= 8'h00;
            16'd783: data <= 8'hF8;
            16'd784: data <= 8'h00;
            16'd785: data <= 8'hF8;
            16'd786: data <= 8'h00;
            16'd787: data <= 8'hF8;
            16'd788: data <= 8'h00;
            16'd789: data <= 8'hF8;
            16'd790: data <= 8'h00;
            16'd791: data <= 8'hF8;
            16'd792: data <= 8'h00;
            16'd793: data <= 8'hF8;
            16'd794: data <= 8'h00;
            16'd795: data <= 8'hF8;
            16'd796: data <= 8'h00;
            16'd797: data <= 8'hF8;
            16'd798: data <= 8'h00;
            16'd799: data <= 8'hF8;
            16'd800: data <= 8'hFF;
            16'd801: data <= 8'hFF;
            16'd802: data <= 8'h00;
            16'd803: data <= 8'hF8;
            16'd804: data <= 8'h00;
            16'd805: data <= 8'hF8;
            16'd806: data <= 8'h00;
            16'd807: data <= 8'hF8;
            16'd808: data <= 8'h00;
            16'd809: data <= 8'hF8;
            16'd810: data <= 8'h00;
            16'd811: data <= 8'hF8;
            16'd812: data <= 8'h00;
            16'd813: data <= 8'hF8;
            16'd814: data <= 8'h00;
            16'd815: data <= 8'hF8;
            16'd816: data <= 8'h00;
            16'd817: data <= 8'hF8;
            16'd818: data <= 8'h00;
            16'd819: data <= 8'hF8;
            16'd820: data <= 8'h00;
            16'd821: data <= 8'hF8;
            16'd822: data <= 8'h00;
            16'd823: data <= 8'hF8;
            16'd824: data <= 8'h00;
            16'd825: data <= 8'hF8;
            16'd826: data <= 8'h00;
            16'd827: data <= 8'hF8;
            16'd828: data <= 8'h00;
            16'd829: data <= 8'hF8;
            16'd830: data <= 8'h00;
            16'd831: data <= 8'hF8;
            16'd832: data <= 8'h00;
            16'd833: data <= 8'hF8;
            16'd834: data <= 8'h00;
            16'd835: data <= 8'hF8;
            16'd836: data <= 8'h00;
            16'd837: data <= 8'hF8;
            16'd838: data <= 8'h00;
            16'd839: data <= 8'hF8;
            16'd840: data <= 8'hFF;
            16'd841: data <= 8'hFF;
            16'd842: data <= 8'h00;
            16'd843: data <= 8'hF8;
            16'd844: data <= 8'h00;
            16'd845: data <= 8'hF8;
            16'd846: data <= 8'h00;
            16'd847: data <= 8'hF8;
            16'd848: data <= 8'h00;
            16'd849: data <= 8'hF8;
            16'd850: data <= 8'h00;
            16'd851: data <= 8'hF8;
            16'd852: data <= 8'h00;
            16'd853: data <= 8'hF8;
            16'd854: data <= 8'h00;
            16'd855: data <= 8'hF8;
            16'd856: data <= 8'h00;
            16'd857: data <= 8'hF8;
            16'd858: data <= 8'h00;
            16'd859: data <= 8'hF8;
            16'd860: data <= 8'h00;
            16'd861: data <= 8'hF8;
            16'd862: data <= 8'h00;
            16'd863: data <= 8'hF8;
            16'd864: data <= 8'h00;
            16'd865: data <= 8'hF8;
            16'd866: data <= 8'h00;
            16'd867: data <= 8'hF8;
            16'd868: data <= 8'h00;
            16'd869: data <= 8'hF8;
            16'd870: data <= 8'h00;
            16'd871: data <= 8'hF8;
            16'd872: data <= 8'h00;
            16'd873: data <= 8'hF8;
            16'd874: data <= 8'h00;
            16'd875: data <= 8'hF8;
            16'd876: data <= 8'h00;
            16'd877: data <= 8'hF8;
            16'd878: data <= 8'h00;
            16'd879: data <= 8'hF8;
            16'd880: data <= 8'hFF;
            16'd881: data <= 8'hFF;
            16'd882: data <= 8'h00;
            16'd883: data <= 8'hF8;
            16'd884: data <= 8'h00;
            16'd885: data <= 8'hF8;
            16'd886: data <= 8'h00;
            16'd887: data <= 8'hF8;
            16'd888: data <= 8'h00;
            16'd889: data <= 8'hF8;
            16'd890: data <= 8'h00;
            16'd891: data <= 8'hF8;
            16'd892: data <= 8'h00;
            16'd893: data <= 8'hF8;
            16'd894: data <= 8'h00;
            16'd895: data <= 8'hF8;
            16'd896: data <= 8'h00;
            16'd897: data <= 8'hF8;
            16'd898: data <= 8'h00;
            16'd899: data <= 8'hF8;
            16'd900: data <= 8'h00;
            16'd901: data <= 8'hF8;
            16'd902: data <= 8'h00;
            16'd903: data <= 8'hF8;
            16'd904: data <= 8'h00;
            16'd905: data <= 8'hF8;
            16'd906: data <= 8'h00;
            16'd907: data <= 8'hF8;
            16'd908: data <= 8'h00;
            16'd909: data <= 8'hF8;
            16'd910: data <= 8'h00;
            16'd911: data <= 8'hF8;
            16'd912: data <= 8'h00;
            16'd913: data <= 8'hF8;
            16'd914: data <= 8'h00;
            16'd915: data <= 8'hF8;
            16'd916: data <= 8'h00;
            16'd917: data <= 8'hF8;
            16'd918: data <= 8'h00;
            16'd919: data <= 8'hF8;
            16'd920: data <= 8'hFF;
            16'd921: data <= 8'hFF;
            16'd922: data <= 8'h00;
            16'd923: data <= 8'hF8;
            16'd924: data <= 8'h00;
            16'd925: data <= 8'hF8;
            16'd926: data <= 8'h00;
            16'd927: data <= 8'hF8;
            16'd928: data <= 8'h00;
            16'd929: data <= 8'hF8;
            16'd930: data <= 8'h00;
            16'd931: data <= 8'hF8;
            16'd932: data <= 8'h00;
            16'd933: data <= 8'hF8;
            16'd934: data <= 8'h00;
            16'd935: data <= 8'hF8;
            16'd936: data <= 8'h00;
            16'd937: data <= 8'hF8;
            16'd938: data <= 8'h00;
            16'd939: data <= 8'hF8;
            16'd940: data <= 8'h00;
            16'd941: data <= 8'hF8;
            16'd942: data <= 8'h00;
            16'd943: data <= 8'hF8;
            16'd944: data <= 8'h00;
            16'd945: data <= 8'hF8;
            16'd946: data <= 8'h00;
            16'd947: data <= 8'hF8;
            16'd948: data <= 8'h00;
            16'd949: data <= 8'hF8;
            16'd950: data <= 8'h00;
            16'd951: data <= 8'hF8;
            16'd952: data <= 8'h00;
            16'd953: data <= 8'hF8;
            16'd954: data <= 8'h00;
            16'd955: data <= 8'hF8;
            16'd956: data <= 8'h00;
            16'd957: data <= 8'hF8;
            16'd958: data <= 8'h00;
            16'd959: data <= 8'hF8;
            16'd960: data <= 8'hFF;
            16'd961: data <= 8'hFF;
            16'd962: data <= 8'h00;
            16'd963: data <= 8'hF8;
            16'd964: data <= 8'h00;
            16'd965: data <= 8'hF8;
            16'd966: data <= 8'h00;
            16'd967: data <= 8'hF8;
            16'd968: data <= 8'h00;
            16'd969: data <= 8'hF8;
            16'd970: data <= 8'h00;
            16'd971: data <= 8'hF8;
            16'd972: data <= 8'h00;
            16'd973: data <= 8'hF8;
            16'd974: data <= 8'h00;
            16'd975: data <= 8'hF8;
            16'd976: data <= 8'h00;
            16'd977: data <= 8'hF8;
            16'd978: data <= 8'h00;
            16'd979: data <= 8'hF8;
            16'd980: data <= 8'h00;
            16'd981: data <= 8'hF8;
            16'd982: data <= 8'h00;
            16'd983: data <= 8'hF8;
            16'd984: data <= 8'h00;
            16'd985: data <= 8'hF8;
            16'd986: data <= 8'h00;
            16'd987: data <= 8'hF8;
            16'd988: data <= 8'h00;
            16'd989: data <= 8'hF8;
            16'd990: data <= 8'h00;
            16'd991: data <= 8'hF8;
            16'd992: data <= 8'h00;
            16'd993: data <= 8'hF8;
            16'd994: data <= 8'h00;
            16'd995: data <= 8'hF8;
            16'd996: data <= 8'h00;
            16'd997: data <= 8'hF8;
            16'd998: data <= 8'h00;
            16'd999: data <= 8'hF8;
            16'd1000: data <= 8'hFF;
            16'd1001: data <= 8'hFF;
            16'd1002: data <= 8'h00;
            16'd1003: data <= 8'hF8;
            16'd1004: data <= 8'h00;
            16'd1005: data <= 8'hF8;
            16'd1006: data <= 8'h00;
            16'd1007: data <= 8'hF8;
            16'd1008: data <= 8'h00;
            16'd1009: data <= 8'hF8;
            16'd1010: data <= 8'h00;
            16'd1011: data <= 8'hF8;
            16'd1012: data <= 8'h00;
            16'd1013: data <= 8'hF8;
            16'd1014: data <= 8'h00;
            16'd1015: data <= 8'hF8;
            16'd1016: data <= 8'h00;
            16'd1017: data <= 8'hF8;
            16'd1018: data <= 8'h00;
            16'd1019: data <= 8'hF8;
            16'd1020: data <= 8'h00;
            16'd1021: data <= 8'hF8;
            16'd1022: data <= 8'h00;
            16'd1023: data <= 8'hF8;
            16'd1024: data <= 8'h00;
            16'd1025: data <= 8'hF8;
            16'd1026: data <= 8'h00;
            16'd1027: data <= 8'hF8;
            16'd1028: data <= 8'h00;
            16'd1029: data <= 8'hF8;
            16'd1030: data <= 8'h00;
            16'd1031: data <= 8'hF8;
            16'd1032: data <= 8'h00;
            16'd1033: data <= 8'hF8;
            16'd1034: data <= 8'h00;
            16'd1035: data <= 8'hF8;
            16'd1036: data <= 8'h00;
            16'd1037: data <= 8'hF8;
            16'd1038: data <= 8'h00;
            16'd1039: data <= 8'hF8;
            16'd1040: data <= 8'hFF;
            16'd1041: data <= 8'hFF;
            16'd1042: data <= 8'h00;
            16'd1043: data <= 8'hF8;
            16'd1044: data <= 8'h00;
            16'd1045: data <= 8'hF8;
            16'd1046: data <= 8'h00;
            16'd1047: data <= 8'hF8;
            16'd1048: data <= 8'h00;
            16'd1049: data <= 8'hF8;
            16'd1050: data <= 8'h00;
            16'd1051: data <= 8'hF8;
            16'd1052: data <= 8'h00;
            16'd1053: data <= 8'hF8;
            16'd1054: data <= 8'h00;
            16'd1055: data <= 8'hF8;
            16'd1056: data <= 8'h00;
            16'd1057: data <= 8'hF8;
            16'd1058: data <= 8'h00;
            16'd1059: data <= 8'hF8;
            16'd1060: data <= 8'h00;
            16'd1061: data <= 8'hF8;
            16'd1062: data <= 8'h00;
            16'd1063: data <= 8'hF8;
            16'd1064: data <= 8'h00;
            16'd1065: data <= 8'hF8;
            16'd1066: data <= 8'h00;
            16'd1067: data <= 8'hF8;
            16'd1068: data <= 8'h00;
            16'd1069: data <= 8'hF8;
            16'd1070: data <= 8'h00;
            16'd1071: data <= 8'hF8;
            16'd1072: data <= 8'h00;
            16'd1073: data <= 8'hF8;
            16'd1074: data <= 8'h00;
            16'd1075: data <= 8'hF8;
            16'd1076: data <= 8'h00;
            16'd1077: data <= 8'hF8;
            16'd1078: data <= 8'h00;
            16'd1079: data <= 8'hF8;
            16'd1080: data <= 8'hFF;
            16'd1081: data <= 8'hFF;
            16'd1082: data <= 8'h00;
            16'd1083: data <= 8'hF8;
            16'd1084: data <= 8'h00;
            16'd1085: data <= 8'hF8;
            16'd1086: data <= 8'h00;
            16'd1087: data <= 8'hF8;
            16'd1088: data <= 8'h00;
            16'd1089: data <= 8'hF8;
            16'd1090: data <= 8'h00;
            16'd1091: data <= 8'hF8;
            16'd1092: data <= 8'h00;
            16'd1093: data <= 8'hF8;
            16'd1094: data <= 8'h00;
            16'd1095: data <= 8'hF8;
            16'd1096: data <= 8'h00;
            16'd1097: data <= 8'hF8;
            16'd1098: data <= 8'h00;
            16'd1099: data <= 8'hF8;
            16'd1100: data <= 8'h00;
            16'd1101: data <= 8'hF8;
            16'd1102: data <= 8'h00;
            16'd1103: data <= 8'hF8;
            16'd1104: data <= 8'h00;
            16'd1105: data <= 8'hF8;
            16'd1106: data <= 8'h00;
            16'd1107: data <= 8'hF8;
            16'd1108: data <= 8'h00;
            16'd1109: data <= 8'hF8;
            16'd1110: data <= 8'h00;
            16'd1111: data <= 8'hF8;
            16'd1112: data <= 8'h00;
            16'd1113: data <= 8'hF8;
            16'd1114: data <= 8'h00;
            16'd1115: data <= 8'hF8;
            16'd1116: data <= 8'h00;
            16'd1117: data <= 8'hF8;
            16'd1118: data <= 8'h00;
            16'd1119: data <= 8'hF8;
            16'd1120: data <= 8'hFF;
            16'd1121: data <= 8'hFF;
            16'd1122: data <= 8'h00;
            16'd1123: data <= 8'hF8;
            16'd1124: data <= 8'h00;
            16'd1125: data <= 8'hF8;
            16'd1126: data <= 8'h00;
            16'd1127: data <= 8'hF8;
            16'd1128: data <= 8'h00;
            16'd1129: data <= 8'hF8;
            16'd1130: data <= 8'h00;
            16'd1131: data <= 8'hF8;
            16'd1132: data <= 8'h00;
            16'd1133: data <= 8'hF8;
            16'd1134: data <= 8'h00;
            16'd1135: data <= 8'hF8;
            16'd1136: data <= 8'h00;
            16'd1137: data <= 8'hF8;
            16'd1138: data <= 8'h00;
            16'd1139: data <= 8'hF8;
            16'd1140: data <= 8'h00;
            16'd1141: data <= 8'hF8;
            16'd1142: data <= 8'h00;
            16'd1143: data <= 8'hF8;
            16'd1144: data <= 8'h00;
            16'd1145: data <= 8'hF8;
            16'd1146: data <= 8'h00;
            16'd1147: data <= 8'hF8;
            16'd1148: data <= 8'h00;
            16'd1149: data <= 8'hF8;
            16'd1150: data <= 8'h00;
            16'd1151: data <= 8'hF8;
            16'd1152: data <= 8'h00;
            16'd1153: data <= 8'hF8;
            16'd1154: data <= 8'h00;
            16'd1155: data <= 8'hF8;
            16'd1156: data <= 8'h00;
            16'd1157: data <= 8'hF8;
            16'd1158: data <= 8'h00;
            16'd1159: data <= 8'hF8;
            16'd1160: data <= 8'hFF;
            16'd1161: data <= 8'hFF;
            16'd1162: data <= 8'h00;
            16'd1163: data <= 8'hF8;
            16'd1164: data <= 8'h00;
            16'd1165: data <= 8'hF8;
            16'd1166: data <= 8'h00;
            16'd1167: data <= 8'hF8;
            16'd1168: data <= 8'h00;
            16'd1169: data <= 8'hF8;
            16'd1170: data <= 8'h00;
            16'd1171: data <= 8'hF8;
            16'd1172: data <= 8'h00;
            16'd1173: data <= 8'hF8;
            16'd1174: data <= 8'h00;
            16'd1175: data <= 8'hF8;
            16'd1176: data <= 8'h00;
            16'd1177: data <= 8'hF8;
            16'd1178: data <= 8'h00;
            16'd1179: data <= 8'hF8;
            16'd1180: data <= 8'h00;
            16'd1181: data <= 8'hF8;
            16'd1182: data <= 8'h00;
            16'd1183: data <= 8'hF8;
            16'd1184: data <= 8'h00;
            16'd1185: data <= 8'hF8;
            16'd1186: data <= 8'h00;
            16'd1187: data <= 8'hF8;
            16'd1188: data <= 8'h00;
            16'd1189: data <= 8'hF8;
            16'd1190: data <= 8'h00;
            16'd1191: data <= 8'hF8;
            16'd1192: data <= 8'h00;
            16'd1193: data <= 8'hF8;
            16'd1194: data <= 8'h00;
            16'd1195: data <= 8'hF8;
            16'd1196: data <= 8'h00;
            16'd1197: data <= 8'hF8;
            16'd1198: data <= 8'h00;
            16'd1199: data <= 8'hF8;
            16'd1200: data <= 8'hFF;
            16'd1201: data <= 8'hFF;
            16'd1202: data <= 8'h00;
            16'd1203: data <= 8'hF8;
            16'd1204: data <= 8'h00;
            16'd1205: data <= 8'hF8;
            16'd1206: data <= 8'h00;
            16'd1207: data <= 8'hF8;
            16'd1208: data <= 8'h00;
            16'd1209: data <= 8'hF8;
            16'd1210: data <= 8'h00;
            16'd1211: data <= 8'hF8;
            16'd1212: data <= 8'h00;
            16'd1213: data <= 8'hF8;
            16'd1214: data <= 8'h00;
            16'd1215: data <= 8'hF8;
            16'd1216: data <= 8'h00;
            16'd1217: data <= 8'hF8;
            16'd1218: data <= 8'h00;
            16'd1219: data <= 8'hF8;
            16'd1220: data <= 8'h00;
            16'd1221: data <= 8'hF8;
            16'd1222: data <= 8'h00;
            16'd1223: data <= 8'hF8;
            16'd1224: data <= 8'h00;
            16'd1225: data <= 8'hF8;
            16'd1226: data <= 8'h00;
            16'd1227: data <= 8'hF8;
            16'd1228: data <= 8'h00;
            16'd1229: data <= 8'hF8;
            16'd1230: data <= 8'h00;
            16'd1231: data <= 8'hF8;
            16'd1232: data <= 8'h00;
            16'd1233: data <= 8'hF8;
            16'd1234: data <= 8'h00;
            16'd1235: data <= 8'hF8;
            16'd1236: data <= 8'h00;
            16'd1237: data <= 8'hF8;
            16'd1238: data <= 8'h00;
            16'd1239: data <= 8'hF8;
            16'd1240: data <= 8'hFF;
            16'd1241: data <= 8'hFF;
            16'd1242: data <= 8'h00;
            16'd1243: data <= 8'hF8;
            16'd1244: data <= 8'h00;
            16'd1245: data <= 8'hF8;
            16'd1246: data <= 8'h00;
            16'd1247: data <= 8'hF8;
            16'd1248: data <= 8'h00;
            16'd1249: data <= 8'hF8;
            16'd1250: data <= 8'h00;
            16'd1251: data <= 8'hF8;
            16'd1252: data <= 8'h00;
            16'd1253: data <= 8'hF8;
            16'd1254: data <= 8'h00;
            16'd1255: data <= 8'hF8;
            16'd1256: data <= 8'h00;
            16'd1257: data <= 8'hF8;
            16'd1258: data <= 8'h00;
            16'd1259: data <= 8'hF8;
            16'd1260: data <= 8'h00;
            16'd1261: data <= 8'hF8;
            16'd1262: data <= 8'h00;
            16'd1263: data <= 8'hF8;
            16'd1264: data <= 8'h00;
            16'd1265: data <= 8'hF8;
            16'd1266: data <= 8'h00;
            16'd1267: data <= 8'hF8;
            16'd1268: data <= 8'h00;
            16'd1269: data <= 8'hF8;
            16'd1270: data <= 8'h00;
            16'd1271: data <= 8'hF8;
            16'd1272: data <= 8'h00;
            16'd1273: data <= 8'hF8;
            16'd1274: data <= 8'h00;
            16'd1275: data <= 8'hF8;
            16'd1276: data <= 8'h00;
            16'd1277: data <= 8'hF8;
            16'd1278: data <= 8'h00;
            16'd1279: data <= 8'hF8;
            16'd1280: data <= 8'hFF;
            16'd1281: data <= 8'hFF;
            16'd1282: data <= 8'h00;
            16'd1283: data <= 8'hF8;
            16'd1284: data <= 8'h00;
            16'd1285: data <= 8'hF8;
            16'd1286: data <= 8'h00;
            16'd1287: data <= 8'hF8;
            16'd1288: data <= 8'h00;
            16'd1289: data <= 8'hF8;
            16'd1290: data <= 8'h00;
            16'd1291: data <= 8'hF8;
            16'd1292: data <= 8'h00;
            16'd1293: data <= 8'hF8;
            16'd1294: data <= 8'h00;
            16'd1295: data <= 8'hF8;
            16'd1296: data <= 8'h00;
            16'd1297: data <= 8'hF8;
            16'd1298: data <= 8'h00;
            16'd1299: data <= 8'hF8;
            16'd1300: data <= 8'h00;
            16'd1301: data <= 8'hF8;
            16'd1302: data <= 8'h00;
            16'd1303: data <= 8'hF8;
            16'd1304: data <= 8'h00;
            16'd1305: data <= 8'hF8;
            16'd1306: data <= 8'h00;
            16'd1307: data <= 8'hF8;
            16'd1308: data <= 8'h00;
            16'd1309: data <= 8'hF8;
            16'd1310: data <= 8'h00;
            16'd1311: data <= 8'hF8;
            16'd1312: data <= 8'h00;
            16'd1313: data <= 8'hF8;
            16'd1314: data <= 8'h00;
            16'd1315: data <= 8'hF8;
            16'd1316: data <= 8'h00;
            16'd1317: data <= 8'hF8;
            16'd1318: data <= 8'h00;
            16'd1319: data <= 8'hF8;
            16'd1320: data <= 8'hFF;
            16'd1321: data <= 8'hFF;
            16'd1322: data <= 8'h00;
            16'd1323: data <= 8'hF8;
            16'd1324: data <= 8'h00;
            16'd1325: data <= 8'hF8;
            16'd1326: data <= 8'h00;
            16'd1327: data <= 8'hF8;
            16'd1328: data <= 8'h00;
            16'd1329: data <= 8'hF8;
            16'd1330: data <= 8'h00;
            16'd1331: data <= 8'hF8;
            16'd1332: data <= 8'h00;
            16'd1333: data <= 8'hF8;
            16'd1334: data <= 8'h00;
            16'd1335: data <= 8'hF8;
            16'd1336: data <= 8'h00;
            16'd1337: data <= 8'hF8;
            16'd1338: data <= 8'h00;
            16'd1339: data <= 8'hF8;
            16'd1340: data <= 8'h00;
            16'd1341: data <= 8'hF8;
            16'd1342: data <= 8'h00;
            16'd1343: data <= 8'hF8;
            16'd1344: data <= 8'h00;
            16'd1345: data <= 8'hF8;
            16'd1346: data <= 8'h00;
            16'd1347: data <= 8'hF8;
            16'd1348: data <= 8'h00;
            16'd1349: data <= 8'hF8;
            16'd1350: data <= 8'h00;
            16'd1351: data <= 8'hF8;
            16'd1352: data <= 8'h00;
            16'd1353: data <= 8'hF8;
            16'd1354: data <= 8'h00;
            16'd1355: data <= 8'hF8;
            16'd1356: data <= 8'h00;
            16'd1357: data <= 8'hF8;
            16'd1358: data <= 8'h00;
            16'd1359: data <= 8'hF8;
            16'd1360: data <= 8'hFF;
            16'd1361: data <= 8'hFF;
            16'd1362: data <= 8'h00;
            16'd1363: data <= 8'hF8;
            16'd1364: data <= 8'h00;
            16'd1365: data <= 8'hF8;
            16'd1366: data <= 8'h00;
            16'd1367: data <= 8'hF8;
            16'd1368: data <= 8'h00;
            16'd1369: data <= 8'hF8;
            16'd1370: data <= 8'h00;
            16'd1371: data <= 8'hF8;
            16'd1372: data <= 8'h00;
            16'd1373: data <= 8'hF8;
            16'd1374: data <= 8'h00;
            16'd1375: data <= 8'hF8;
            16'd1376: data <= 8'h00;
            16'd1377: data <= 8'hF8;
            16'd1378: data <= 8'h00;
            16'd1379: data <= 8'hF8;
            16'd1380: data <= 8'h00;
            16'd1381: data <= 8'hF8;
            16'd1382: data <= 8'h00;
            16'd1383: data <= 8'hF8;
            16'd1384: data <= 8'h00;
            16'd1385: data <= 8'hF8;
            16'd1386: data <= 8'h00;
            16'd1387: data <= 8'hF8;
            16'd1388: data <= 8'h00;
            16'd1389: data <= 8'hF8;
            16'd1390: data <= 8'h00;
            16'd1391: data <= 8'hF8;
            16'd1392: data <= 8'h00;
            16'd1393: data <= 8'hF8;
            16'd1394: data <= 8'h00;
            16'd1395: data <= 8'hF8;
            16'd1396: data <= 8'h00;
            16'd1397: data <= 8'hF8;
            16'd1398: data <= 8'h00;
            16'd1399: data <= 8'hF8;
            16'd1400: data <= 8'hFF;
            16'd1401: data <= 8'hFF;
            16'd1402: data <= 8'h00;
            16'd1403: data <= 8'hF8;
            16'd1404: data <= 8'h00;
            16'd1405: data <= 8'hF8;
            16'd1406: data <= 8'h00;
            16'd1407: data <= 8'hF8;
            16'd1408: data <= 8'h00;
            16'd1409: data <= 8'hF8;
            16'd1410: data <= 8'h00;
            16'd1411: data <= 8'hF8;
            16'd1412: data <= 8'h00;
            16'd1413: data <= 8'hF8;
            16'd1414: data <= 8'h00;
            16'd1415: data <= 8'hF8;
            16'd1416: data <= 8'h00;
            16'd1417: data <= 8'hF8;
            16'd1418: data <= 8'h00;
            16'd1419: data <= 8'hF8;
            16'd1420: data <= 8'h00;
            16'd1421: data <= 8'hF8;
            16'd1422: data <= 8'h00;
            16'd1423: data <= 8'hF8;
            16'd1424: data <= 8'h00;
            16'd1425: data <= 8'hF8;
            16'd1426: data <= 8'h00;
            16'd1427: data <= 8'hF8;
            16'd1428: data <= 8'h00;
            16'd1429: data <= 8'hF8;
            16'd1430: data <= 8'h00;
            16'd1431: data <= 8'hF8;
            16'd1432: data <= 8'h00;
            16'd1433: data <= 8'hF8;
            16'd1434: data <= 8'h00;
            16'd1435: data <= 8'hF8;
            16'd1436: data <= 8'h00;
            16'd1437: data <= 8'hF8;
            16'd1438: data <= 8'h00;
            16'd1439: data <= 8'hF8;
            16'd1440: data <= 8'hFF;
            16'd1441: data <= 8'hFF;
            16'd1442: data <= 8'h00;
            16'd1443: data <= 8'hF8;
            16'd1444: data <= 8'h00;
            16'd1445: data <= 8'hF8;
            16'd1446: data <= 8'h00;
            16'd1447: data <= 8'hF8;
            16'd1448: data <= 8'h00;
            16'd1449: data <= 8'hF8;
            16'd1450: data <= 8'h00;
            16'd1451: data <= 8'hF8;
            16'd1452: data <= 8'h00;
            16'd1453: data <= 8'hF8;
            16'd1454: data <= 8'h00;
            16'd1455: data <= 8'hF8;
            16'd1456: data <= 8'h00;
            16'd1457: data <= 8'hF8;
            16'd1458: data <= 8'h00;
            16'd1459: data <= 8'hF8;
            16'd1460: data <= 8'h00;
            16'd1461: data <= 8'hF8;
            16'd1462: data <= 8'h00;
            16'd1463: data <= 8'hF8;
            16'd1464: data <= 8'h00;
            16'd1465: data <= 8'hF8;
            16'd1466: data <= 8'h00;
            16'd1467: data <= 8'hF8;
            16'd1468: data <= 8'h00;
            16'd1469: data <= 8'hF8;
            16'd1470: data <= 8'h00;
            16'd1471: data <= 8'hF8;
            16'd1472: data <= 8'h00;
            16'd1473: data <= 8'hF8;
            16'd1474: data <= 8'h00;
            16'd1475: data <= 8'hF8;
            16'd1476: data <= 8'h00;
            16'd1477: data <= 8'hF8;
            16'd1478: data <= 8'h00;
            16'd1479: data <= 8'hF8;
            16'd1480: data <= 8'hFF;
            16'd1481: data <= 8'hFF;
            16'd1482: data <= 8'h00;
            16'd1483: data <= 8'hF8;
            16'd1484: data <= 8'h00;
            16'd1485: data <= 8'hF8;
            16'd1486: data <= 8'h00;
            16'd1487: data <= 8'hF8;
            16'd1488: data <= 8'h00;
            16'd1489: data <= 8'hF8;
            16'd1490: data <= 8'h00;
            16'd1491: data <= 8'hF8;
            16'd1492: data <= 8'h00;
            16'd1493: data <= 8'hF8;
            16'd1494: data <= 8'h00;
            16'd1495: data <= 8'hF8;
            16'd1496: data <= 8'h00;
            16'd1497: data <= 8'hF8;
            16'd1498: data <= 8'h00;
            16'd1499: data <= 8'hF8;
            16'd1500: data <= 8'h00;
            16'd1501: data <= 8'hF8;
            16'd1502: data <= 8'h00;
            16'd1503: data <= 8'hF8;
            16'd1504: data <= 8'h00;
            16'd1505: data <= 8'hF8;
            16'd1506: data <= 8'h00;
            16'd1507: data <= 8'hF8;
            16'd1508: data <= 8'h00;
            16'd1509: data <= 8'hF8;
            16'd1510: data <= 8'h00;
            16'd1511: data <= 8'hF8;
            16'd1512: data <= 8'h00;
            16'd1513: data <= 8'hF8;
            16'd1514: data <= 8'h00;
            16'd1515: data <= 8'hF8;
            16'd1516: data <= 8'h00;
            16'd1517: data <= 8'hF8;
            16'd1518: data <= 8'h00;
            16'd1519: data <= 8'hF8;
            16'd1520: data <= 8'hFF;
            16'd1521: data <= 8'hFF;
            16'd1522: data <= 8'h00;
            16'd1523: data <= 8'hF8;
            16'd1524: data <= 8'h00;
            16'd1525: data <= 8'hF8;
            16'd1526: data <= 8'h00;
            16'd1527: data <= 8'hF8;
            16'd1528: data <= 8'h00;
            16'd1529: data <= 8'hF8;
            16'd1530: data <= 8'h00;
            16'd1531: data <= 8'hF8;
            16'd1532: data <= 8'h00;
            16'd1533: data <= 8'hF8;
            16'd1534: data <= 8'h00;
            16'd1535: data <= 8'hF8;
            16'd1536: data <= 8'h00;
            16'd1537: data <= 8'hF8;
            16'd1538: data <= 8'h00;
            16'd1539: data <= 8'hF8;
            16'd1540: data <= 8'h00;
            16'd1541: data <= 8'hF8;
            16'd1542: data <= 8'h00;
            16'd1543: data <= 8'hF8;
            16'd1544: data <= 8'h00;
            16'd1545: data <= 8'hF8;
            16'd1546: data <= 8'h00;
            16'd1547: data <= 8'hF8;
            16'd1548: data <= 8'h00;
            16'd1549: data <= 8'hF8;
            16'd1550: data <= 8'h00;
            16'd1551: data <= 8'hF8;
            16'd1552: data <= 8'h00;
            16'd1553: data <= 8'hF8;
            16'd1554: data <= 8'h00;
            16'd1555: data <= 8'hF8;
            16'd1556: data <= 8'h00;
            16'd1557: data <= 8'hF8;
            16'd1558: data <= 8'h00;
            16'd1559: data <= 8'hF8;
            16'd1560: data <= 8'hFF;
            16'd1561: data <= 8'hFF;
            16'd1562: data <= 8'h00;
            16'd1563: data <= 8'hF8;
            16'd1564: data <= 8'h00;
            16'd1565: data <= 8'hF8;
            16'd1566: data <= 8'h00;
            16'd1567: data <= 8'hF8;
            16'd1568: data <= 8'h00;
            16'd1569: data <= 8'hF8;
            16'd1570: data <= 8'h00;
            16'd1571: data <= 8'hF8;
            16'd1572: data <= 8'h00;
            16'd1573: data <= 8'hF8;
            16'd1574: data <= 8'h00;
            16'd1575: data <= 8'hF8;
            16'd1576: data <= 8'h00;
            16'd1577: data <= 8'hF8;
            16'd1578: data <= 8'h00;
            16'd1579: data <= 8'hF8;
            16'd1580: data <= 8'h00;
            16'd1581: data <= 8'hF8;
            16'd1582: data <= 8'h00;
            16'd1583: data <= 8'hF8;
            16'd1584: data <= 8'h00;
            16'd1585: data <= 8'hF8;
            16'd1586: data <= 8'h00;
            16'd1587: data <= 8'hF8;
            16'd1588: data <= 8'h00;
            16'd1589: data <= 8'hF8;
            16'd1590: data <= 8'h00;
            16'd1591: data <= 8'hF8;
            16'd1592: data <= 8'h00;
            16'd1593: data <= 8'hF8;
            16'd1594: data <= 8'h00;
            16'd1595: data <= 8'hF8;
            16'd1596: data <= 8'h00;
            16'd1597: data <= 8'hF8;
            16'd1598: data <= 8'h00;
            16'd1599: data <= 8'hF8;
            16'd1600: data <= 8'hFF;
            16'd1601: data <= 8'hFF;
            16'd1602: data <= 8'h00;
            16'd1603: data <= 8'hF8;
            16'd1604: data <= 8'h00;
            16'd1605: data <= 8'hF8;
            16'd1606: data <= 8'h00;
            16'd1607: data <= 8'hF8;
            16'd1608: data <= 8'h00;
            16'd1609: data <= 8'hF8;
            16'd1610: data <= 8'h00;
            16'd1611: data <= 8'hF8;
            16'd1612: data <= 8'h00;
            16'd1613: data <= 8'hF8;
            16'd1614: data <= 8'h00;
            16'd1615: data <= 8'hF8;
            16'd1616: data <= 8'h00;
            16'd1617: data <= 8'hF8;
            16'd1618: data <= 8'h00;
            16'd1619: data <= 8'hF8;
            16'd1620: data <= 8'h00;
            16'd1621: data <= 8'hF8;
            16'd1622: data <= 8'h00;
            16'd1623: data <= 8'hF8;
            16'd1624: data <= 8'h00;
            16'd1625: data <= 8'hF8;
            16'd1626: data <= 8'h00;
            16'd1627: data <= 8'hF8;
            16'd1628: data <= 8'h00;
            16'd1629: data <= 8'hF8;
            16'd1630: data <= 8'h00;
            16'd1631: data <= 8'hF8;
            16'd1632: data <= 8'h00;
            16'd1633: data <= 8'hF8;
            16'd1634: data <= 8'h00;
            16'd1635: data <= 8'hF8;
            16'd1636: data <= 8'h00;
            16'd1637: data <= 8'hF8;
            16'd1638: data <= 8'h00;
            16'd1639: data <= 8'hF8;
            16'd1640: data <= 8'hFF;
            16'd1641: data <= 8'hFF;
            16'd1642: data <= 8'h00;
            16'd1643: data <= 8'hF8;
            16'd1644: data <= 8'h00;
            16'd1645: data <= 8'hF8;
            16'd1646: data <= 8'h00;
            16'd1647: data <= 8'hF8;
            16'd1648: data <= 8'h00;
            16'd1649: data <= 8'hF8;
            16'd1650: data <= 8'h00;
            16'd1651: data <= 8'hF8;
            16'd1652: data <= 8'h00;
            16'd1653: data <= 8'hF8;
            16'd1654: data <= 8'h00;
            16'd1655: data <= 8'hF8;
            16'd1656: data <= 8'h00;
            16'd1657: data <= 8'hF8;
            16'd1658: data <= 8'h00;
            16'd1659: data <= 8'hF8;
            16'd1660: data <= 8'h00;
            16'd1661: data <= 8'hF8;
            16'd1662: data <= 8'h00;
            16'd1663: data <= 8'hF8;
            16'd1664: data <= 8'h00;
            16'd1665: data <= 8'hF8;
            16'd1666: data <= 8'h00;
            16'd1667: data <= 8'hF8;
            16'd1668: data <= 8'h00;
            16'd1669: data <= 8'hF8;
            16'd1670: data <= 8'h00;
            16'd1671: data <= 8'hF8;
            16'd1672: data <= 8'h00;
            16'd1673: data <= 8'hF8;
            16'd1674: data <= 8'h00;
            16'd1675: data <= 8'hF8;
            16'd1676: data <= 8'h00;
            16'd1677: data <= 8'hF8;
            16'd1678: data <= 8'h00;
            16'd1679: data <= 8'hF8;
            16'd1680: data <= 8'hFF;
            16'd1681: data <= 8'hFF;
            16'd1682: data <= 8'h00;
            16'd1683: data <= 8'hF8;
            16'd1684: data <= 8'h00;
            16'd1685: data <= 8'hF8;
            16'd1686: data <= 8'h00;
            16'd1687: data <= 8'hF8;
            16'd1688: data <= 8'h00;
            16'd1689: data <= 8'hF8;
            16'd1690: data <= 8'h00;
            16'd1691: data <= 8'hF8;
            16'd1692: data <= 8'h00;
            16'd1693: data <= 8'hF8;
            16'd1694: data <= 8'h00;
            16'd1695: data <= 8'hF8;
            16'd1696: data <= 8'h00;
            16'd1697: data <= 8'hF8;
            16'd1698: data <= 8'h00;
            16'd1699: data <= 8'hF8;
            16'd1700: data <= 8'h00;
            16'd1701: data <= 8'hF8;
            16'd1702: data <= 8'h00;
            16'd1703: data <= 8'hF8;
            16'd1704: data <= 8'h00;
            16'd1705: data <= 8'hF8;
            16'd1706: data <= 8'h00;
            16'd1707: data <= 8'hF8;
            16'd1708: data <= 8'h00;
            16'd1709: data <= 8'hF8;
            16'd1710: data <= 8'h00;
            16'd1711: data <= 8'hF8;
            16'd1712: data <= 8'h00;
            16'd1713: data <= 8'hF8;
            16'd1714: data <= 8'h00;
            16'd1715: data <= 8'hF8;
            16'd1716: data <= 8'h00;
            16'd1717: data <= 8'hF8;
            16'd1718: data <= 8'h00;
            16'd1719: data <= 8'hF8;
            16'd1720: data <= 8'hFF;
            16'd1721: data <= 8'hFF;
            16'd1722: data <= 8'h00;
            16'd1723: data <= 8'hF8;
            16'd1724: data <= 8'h00;
            16'd1725: data <= 8'hF8;
            16'd1726: data <= 8'h00;
            16'd1727: data <= 8'hF8;
            16'd1728: data <= 8'h00;
            16'd1729: data <= 8'hF8;
            16'd1730: data <= 8'h00;
            16'd1731: data <= 8'hF8;
            16'd1732: data <= 8'h00;
            16'd1733: data <= 8'hF8;
            16'd1734: data <= 8'h00;
            16'd1735: data <= 8'hF8;
            16'd1736: data <= 8'h00;
            16'd1737: data <= 8'hF8;
            16'd1738: data <= 8'h00;
            16'd1739: data <= 8'hF8;
            16'd1740: data <= 8'h00;
            16'd1741: data <= 8'hF8;
            16'd1742: data <= 8'h00;
            16'd1743: data <= 8'hF8;
            16'd1744: data <= 8'h00;
            16'd1745: data <= 8'hF8;
            16'd1746: data <= 8'h00;
            16'd1747: data <= 8'hF8;
            16'd1748: data <= 8'h00;
            16'd1749: data <= 8'hF8;
            16'd1750: data <= 8'h00;
            16'd1751: data <= 8'hF8;
            16'd1752: data <= 8'h00;
            16'd1753: data <= 8'hF8;
            16'd1754: data <= 8'h00;
            16'd1755: data <= 8'hF8;
            16'd1756: data <= 8'h00;
            16'd1757: data <= 8'hF8;
            16'd1758: data <= 8'h00;
            16'd1759: data <= 8'hF8;
            16'd1760: data <= 8'hFF;
            16'd1761: data <= 8'hFF;
            16'd1762: data <= 8'h00;
            16'd1763: data <= 8'hF8;
            16'd1764: data <= 8'h00;
            16'd1765: data <= 8'hF8;
            16'd1766: data <= 8'h00;
            16'd1767: data <= 8'hF8;
            16'd1768: data <= 8'h00;
            16'd1769: data <= 8'hF8;
            16'd1770: data <= 8'h00;
            16'd1771: data <= 8'hF8;
            16'd1772: data <= 8'h00;
            16'd1773: data <= 8'hF8;
            16'd1774: data <= 8'h00;
            16'd1775: data <= 8'hF8;
            16'd1776: data <= 8'h00;
            16'd1777: data <= 8'hF8;
            16'd1778: data <= 8'h00;
            16'd1779: data <= 8'hF8;
            16'd1780: data <= 8'h00;
            16'd1781: data <= 8'hF8;
            16'd1782: data <= 8'h00;
            16'd1783: data <= 8'hF8;
            16'd1784: data <= 8'h00;
            16'd1785: data <= 8'hF8;
            16'd1786: data <= 8'h00;
            16'd1787: data <= 8'hF8;
            16'd1788: data <= 8'h00;
            16'd1789: data <= 8'hF8;
            16'd1790: data <= 8'h00;
            16'd1791: data <= 8'hF8;
            16'd1792: data <= 8'h00;
            16'd1793: data <= 8'hF8;
            16'd1794: data <= 8'h00;
            16'd1795: data <= 8'hF8;
            16'd1796: data <= 8'h00;
            16'd1797: data <= 8'hF8;
            16'd1798: data <= 8'h00;
            16'd1799: data <= 8'hF8;
            16'd1800: data <= 8'hFF;
            16'd1801: data <= 8'hFF;
            16'd1802: data <= 8'h00;
            16'd1803: data <= 8'hF8;
            16'd1804: data <= 8'h00;
            16'd1805: data <= 8'hF8;
            16'd1806: data <= 8'h00;
            16'd1807: data <= 8'hF8;
            16'd1808: data <= 8'h00;
            16'd1809: data <= 8'hF8;
            16'd1810: data <= 8'h00;
            16'd1811: data <= 8'hF8;
            16'd1812: data <= 8'h00;
            16'd1813: data <= 8'hF8;
            16'd1814: data <= 8'h00;
            16'd1815: data <= 8'hF8;
            16'd1816: data <= 8'h00;
            16'd1817: data <= 8'hF8;
            16'd1818: data <= 8'h00;
            16'd1819: data <= 8'hF8;
            16'd1820: data <= 8'h00;
            16'd1821: data <= 8'hF8;
            16'd1822: data <= 8'h00;
            16'd1823: data <= 8'hF8;
            16'd1824: data <= 8'h00;
            16'd1825: data <= 8'hF8;
            16'd1826: data <= 8'h00;
            16'd1827: data <= 8'hF8;
            16'd1828: data <= 8'h00;
            16'd1829: data <= 8'hF8;
            16'd1830: data <= 8'h00;
            16'd1831: data <= 8'hF8;
            16'd1832: data <= 8'h00;
            16'd1833: data <= 8'hF8;
            16'd1834: data <= 8'h00;
            16'd1835: data <= 8'hF8;
            16'd1836: data <= 8'h00;
            16'd1837: data <= 8'hF8;
            16'd1838: data <= 8'h00;
            16'd1839: data <= 8'hF8;
            16'd1840: data <= 8'hFF;
            16'd1841: data <= 8'hFF;
            16'd1842: data <= 8'h00;
            16'd1843: data <= 8'hF8;
            16'd1844: data <= 8'h00;
            16'd1845: data <= 8'hF8;
            16'd1846: data <= 8'h00;
            16'd1847: data <= 8'hF8;
            16'd1848: data <= 8'h00;
            16'd1849: data <= 8'hF8;
            16'd1850: data <= 8'h00;
            16'd1851: data <= 8'hF8;
            16'd1852: data <= 8'h00;
            16'd1853: data <= 8'hF8;
            16'd1854: data <= 8'h00;
            16'd1855: data <= 8'hF8;
            16'd1856: data <= 8'h00;
            16'd1857: data <= 8'hF8;
            16'd1858: data <= 8'h00;
            16'd1859: data <= 8'hF8;
            16'd1860: data <= 8'h00;
            16'd1861: data <= 8'hF8;
            16'd1862: data <= 8'h00;
            16'd1863: data <= 8'hF8;
            16'd1864: data <= 8'h00;
            16'd1865: data <= 8'hF8;
            16'd1866: data <= 8'h00;
            16'd1867: data <= 8'hF8;
            16'd1868: data <= 8'h00;
            16'd1869: data <= 8'hF8;
            16'd1870: data <= 8'h00;
            16'd1871: data <= 8'hF8;
            16'd1872: data <= 8'h00;
            16'd1873: data <= 8'hF8;
            16'd1874: data <= 8'h00;
            16'd1875: data <= 8'hF8;
            16'd1876: data <= 8'h00;
            16'd1877: data <= 8'hF8;
            16'd1878: data <= 8'h00;
            16'd1879: data <= 8'hF8;
            16'd1880: data <= 8'hFF;
            16'd1881: data <= 8'hFF;
            16'd1882: data <= 8'h00;
            16'd1883: data <= 8'hF8;
            16'd1884: data <= 8'h00;
            16'd1885: data <= 8'hF8;
            16'd1886: data <= 8'h00;
            16'd1887: data <= 8'hF8;
            16'd1888: data <= 8'h00;
            16'd1889: data <= 8'hF8;
            16'd1890: data <= 8'h00;
            16'd1891: data <= 8'hF8;
            16'd1892: data <= 8'h00;
            16'd1893: data <= 8'hF8;
            16'd1894: data <= 8'h00;
            16'd1895: data <= 8'hF8;
            16'd1896: data <= 8'h00;
            16'd1897: data <= 8'hF8;
            16'd1898: data <= 8'h00;
            16'd1899: data <= 8'hF8;
            16'd1900: data <= 8'h00;
            16'd1901: data <= 8'hF8;
            16'd1902: data <= 8'h00;
            16'd1903: data <= 8'hF8;
            16'd1904: data <= 8'h00;
            16'd1905: data <= 8'hF8;
            16'd1906: data <= 8'h00;
            16'd1907: data <= 8'hF8;
            16'd1908: data <= 8'h00;
            16'd1909: data <= 8'hF8;
            16'd1910: data <= 8'h00;
            16'd1911: data <= 8'hF8;
            16'd1912: data <= 8'h00;
            16'd1913: data <= 8'hF8;
            16'd1914: data <= 8'h00;
            16'd1915: data <= 8'hF8;
            16'd1916: data <= 8'h00;
            16'd1917: data <= 8'hF8;
            16'd1918: data <= 8'h00;
            16'd1919: data <= 8'hF8;
            16'd1920: data <= 8'hFF;
            16'd1921: data <= 8'hFF;
            16'd1922: data <= 8'h00;
            16'd1923: data <= 8'hF8;
            16'd1924: data <= 8'h00;
            16'd1925: data <= 8'hF8;
            16'd1926: data <= 8'h00;
            16'd1927: data <= 8'hF8;
            16'd1928: data <= 8'h00;
            16'd1929: data <= 8'hF8;
            16'd1930: data <= 8'h00;
            16'd1931: data <= 8'hF8;
            16'd1932: data <= 8'h00;
            16'd1933: data <= 8'hF8;
            16'd1934: data <= 8'h00;
            16'd1935: data <= 8'hF8;
            16'd1936: data <= 8'h00;
            16'd1937: data <= 8'hF8;
            16'd1938: data <= 8'h00;
            16'd1939: data <= 8'hF8;
            16'd1940: data <= 8'h00;
            16'd1941: data <= 8'hF8;
            16'd1942: data <= 8'h00;
            16'd1943: data <= 8'hF8;
            16'd1944: data <= 8'h00;
            16'd1945: data <= 8'hF8;
            16'd1946: data <= 8'h00;
            16'd1947: data <= 8'hF8;
            16'd1948: data <= 8'h00;
            16'd1949: data <= 8'hF8;
            16'd1950: data <= 8'h00;
            16'd1951: data <= 8'hF8;
            16'd1952: data <= 8'h00;
            16'd1953: data <= 8'hF8;
            16'd1954: data <= 8'h00;
            16'd1955: data <= 8'hF8;
            16'd1956: data <= 8'h00;
            16'd1957: data <= 8'hF8;
            16'd1958: data <= 8'h00;
            16'd1959: data <= 8'hF8;
            16'd1960: data <= 8'hFF;
            16'd1961: data <= 8'hFF;
            16'd1962: data <= 8'h00;
            16'd1963: data <= 8'hF8;
            16'd1964: data <= 8'h00;
            16'd1965: data <= 8'hF8;
            16'd1966: data <= 8'h00;
            16'd1967: data <= 8'hF8;
            16'd1968: data <= 8'h00;
            16'd1969: data <= 8'hF8;
            16'd1970: data <= 8'h00;
            16'd1971: data <= 8'hF8;
            16'd1972: data <= 8'h00;
            16'd1973: data <= 8'hF8;
            16'd1974: data <= 8'h00;
            16'd1975: data <= 8'hF8;
            16'd1976: data <= 8'h00;
            16'd1977: data <= 8'hF8;
            16'd1978: data <= 8'h00;
            16'd1979: data <= 8'hF8;
            16'd1980: data <= 8'h00;
            16'd1981: data <= 8'hF8;
            16'd1982: data <= 8'h00;
            16'd1983: data <= 8'hF8;
            16'd1984: data <= 8'h00;
            16'd1985: data <= 8'hF8;
            16'd1986: data <= 8'h00;
            16'd1987: data <= 8'hF8;
            16'd1988: data <= 8'h00;
            16'd1989: data <= 8'hF8;
            16'd1990: data <= 8'h00;
            16'd1991: data <= 8'hF8;
            16'd1992: data <= 8'h00;
            16'd1993: data <= 8'hF8;
            16'd1994: data <= 8'h00;
            16'd1995: data <= 8'hF8;
            16'd1996: data <= 8'h00;
            16'd1997: data <= 8'hF8;
            16'd1998: data <= 8'h00;
            16'd1999: data <= 8'hF8;
            16'd2000: data <= 8'hFF;
            16'd2001: data <= 8'hFF;
            16'd2002: data <= 8'h00;
            16'd2003: data <= 8'hF8;
            16'd2004: data <= 8'h00;
            16'd2005: data <= 8'hF8;
            16'd2006: data <= 8'h00;
            16'd2007: data <= 8'hF8;
            16'd2008: data <= 8'h00;
            16'd2009: data <= 8'hF8;
            16'd2010: data <= 8'h00;
            16'd2011: data <= 8'hF8;
            16'd2012: data <= 8'h00;
            16'd2013: data <= 8'hF8;
            16'd2014: data <= 8'h00;
            16'd2015: data <= 8'hF8;
            16'd2016: data <= 8'h00;
            16'd2017: data <= 8'hF8;
            16'd2018: data <= 8'h00;
            16'd2019: data <= 8'hF8;
            16'd2020: data <= 8'h00;
            16'd2021: data <= 8'hF8;
            16'd2022: data <= 8'h00;
            16'd2023: data <= 8'hF8;
            16'd2024: data <= 8'h00;
            16'd2025: data <= 8'hF8;
            16'd2026: data <= 8'h00;
            16'd2027: data <= 8'hF8;
            16'd2028: data <= 8'h00;
            16'd2029: data <= 8'hF8;
            16'd2030: data <= 8'h00;
            16'd2031: data <= 8'hF8;
            16'd2032: data <= 8'h00;
            16'd2033: data <= 8'hF8;
            16'd2034: data <= 8'h00;
            16'd2035: data <= 8'hF8;
            16'd2036: data <= 8'h00;
            16'd2037: data <= 8'hF8;
            16'd2038: data <= 8'h00;
            16'd2039: data <= 8'hF8;
            16'd2040: data <= 8'hFF;
            16'd2041: data <= 8'hFF;
            16'd2042: data <= 8'h00;
            16'd2043: data <= 8'hF8;
            16'd2044: data <= 8'h00;
            16'd2045: data <= 8'hF8;
            16'd2046: data <= 8'h00;
            16'd2047: data <= 8'hF8;
            16'd2048: data <= 8'h00;
            16'd2049: data <= 8'hF8;
            16'd2050: data <= 8'h00;
            16'd2051: data <= 8'hF8;
            16'd2052: data <= 8'h00;
            16'd2053: data <= 8'hF8;
            16'd2054: data <= 8'h00;
            16'd2055: data <= 8'hF8;
            16'd2056: data <= 8'h00;
            16'd2057: data <= 8'hF8;
            16'd2058: data <= 8'h00;
            16'd2059: data <= 8'hF8;
            16'd2060: data <= 8'h00;
            16'd2061: data <= 8'hF8;
            16'd2062: data <= 8'h00;
            16'd2063: data <= 8'hF8;
            16'd2064: data <= 8'h00;
            16'd2065: data <= 8'hF8;
            16'd2066: data <= 8'h00;
            16'd2067: data <= 8'hF8;
            16'd2068: data <= 8'h00;
            16'd2069: data <= 8'hF8;
            16'd2070: data <= 8'h00;
            16'd2071: data <= 8'hF8;
            16'd2072: data <= 8'h00;
            16'd2073: data <= 8'hF8;
            16'd2074: data <= 8'h00;
            16'd2075: data <= 8'hF8;
            16'd2076: data <= 8'h00;
            16'd2077: data <= 8'hF8;
            16'd2078: data <= 8'h00;
            16'd2079: data <= 8'hF8;
            16'd2080: data <= 8'hFF;
            16'd2081: data <= 8'hFF;
            16'd2082: data <= 8'h00;
            16'd2083: data <= 8'hF8;
            16'd2084: data <= 8'h00;
            16'd2085: data <= 8'hF8;
            16'd2086: data <= 8'h00;
            16'd2087: data <= 8'hF8;
            16'd2088: data <= 8'h00;
            16'd2089: data <= 8'hF8;
            16'd2090: data <= 8'h00;
            16'd2091: data <= 8'hF8;
            16'd2092: data <= 8'h00;
            16'd2093: data <= 8'hF8;
            16'd2094: data <= 8'h00;
            16'd2095: data <= 8'hF8;
            16'd2096: data <= 8'h00;
            16'd2097: data <= 8'hF8;
            16'd2098: data <= 8'h00;
            16'd2099: data <= 8'hF8;
            16'd2100: data <= 8'h00;
            16'd2101: data <= 8'hF8;
            16'd2102: data <= 8'h00;
            16'd2103: data <= 8'hF8;
            16'd2104: data <= 8'h00;
            16'd2105: data <= 8'hF8;
            16'd2106: data <= 8'h00;
            16'd2107: data <= 8'hF8;
            16'd2108: data <= 8'h00;
            16'd2109: data <= 8'hF8;
            16'd2110: data <= 8'h00;
            16'd2111: data <= 8'hF8;
            16'd2112: data <= 8'h00;
            16'd2113: data <= 8'hF8;
            16'd2114: data <= 8'h00;
            16'd2115: data <= 8'hF8;
            16'd2116: data <= 8'h00;
            16'd2117: data <= 8'hF8;
            16'd2118: data <= 8'h00;
            16'd2119: data <= 8'hF8;
            16'd2120: data <= 8'hFF;
            16'd2121: data <= 8'hFF;
            16'd2122: data <= 8'h00;
            16'd2123: data <= 8'hF8;
            16'd2124: data <= 8'h00;
            16'd2125: data <= 8'hF8;
            16'd2126: data <= 8'h00;
            16'd2127: data <= 8'hF8;
            16'd2128: data <= 8'h00;
            16'd2129: data <= 8'hF8;
            16'd2130: data <= 8'h00;
            16'd2131: data <= 8'hF8;
            16'd2132: data <= 8'h00;
            16'd2133: data <= 8'hF8;
            16'd2134: data <= 8'h00;
            16'd2135: data <= 8'hF8;
            16'd2136: data <= 8'h00;
            16'd2137: data <= 8'hF8;
            16'd2138: data <= 8'h00;
            16'd2139: data <= 8'hF8;
            16'd2140: data <= 8'h00;
            16'd2141: data <= 8'hF8;
            16'd2142: data <= 8'h00;
            16'd2143: data <= 8'hF8;
            16'd2144: data <= 8'h00;
            16'd2145: data <= 8'hF8;
            16'd2146: data <= 8'h00;
            16'd2147: data <= 8'hF8;
            16'd2148: data <= 8'h00;
            16'd2149: data <= 8'hF8;
            16'd2150: data <= 8'h00;
            16'd2151: data <= 8'hF8;
            16'd2152: data <= 8'h00;
            16'd2153: data <= 8'hF8;
            16'd2154: data <= 8'h00;
            16'd2155: data <= 8'hF8;
            16'd2156: data <= 8'h00;
            16'd2157: data <= 8'hF8;
            16'd2158: data <= 8'h00;
            16'd2159: data <= 8'hF8;
            16'd2160: data <= 8'hFF;
            16'd2161: data <= 8'hFF;
            16'd2162: data <= 8'h00;
            16'd2163: data <= 8'hF8;
            16'd2164: data <= 8'h00;
            16'd2165: data <= 8'hF8;
            16'd2166: data <= 8'h00;
            16'd2167: data <= 8'hF8;
            16'd2168: data <= 8'h00;
            16'd2169: data <= 8'hF8;
            16'd2170: data <= 8'h00;
            16'd2171: data <= 8'hF8;
            16'd2172: data <= 8'h00;
            16'd2173: data <= 8'hF8;
            16'd2174: data <= 8'h00;
            16'd2175: data <= 8'hF8;
            16'd2176: data <= 8'h00;
            16'd2177: data <= 8'hF8;
            16'd2178: data <= 8'h00;
            16'd2179: data <= 8'hF8;
            16'd2180: data <= 8'h00;
            16'd2181: data <= 8'hF8;
            16'd2182: data <= 8'h00;
            16'd2183: data <= 8'hF8;
            16'd2184: data <= 8'h00;
            16'd2185: data <= 8'hF8;
            16'd2186: data <= 8'h00;
            16'd2187: data <= 8'hF8;
            16'd2188: data <= 8'h00;
            16'd2189: data <= 8'hF8;
            16'd2190: data <= 8'h00;
            16'd2191: data <= 8'hF8;
            16'd2192: data <= 8'h00;
            16'd2193: data <= 8'hF8;
            16'd2194: data <= 8'h00;
            16'd2195: data <= 8'hF8;
            16'd2196: data <= 8'h00;
            16'd2197: data <= 8'hF8;
            16'd2198: data <= 8'h00;
            16'd2199: data <= 8'hF8;
            16'd2200: data <= 8'hFF;
            16'd2201: data <= 8'hFF;
            16'd2202: data <= 8'h00;
            16'd2203: data <= 8'hF8;
            16'd2204: data <= 8'h00;
            16'd2205: data <= 8'hF8;
            16'd2206: data <= 8'h00;
            16'd2207: data <= 8'hF8;
            16'd2208: data <= 8'h00;
            16'd2209: data <= 8'hF8;
            16'd2210: data <= 8'h00;
            16'd2211: data <= 8'hF8;
            16'd2212: data <= 8'h00;
            16'd2213: data <= 8'hF8;
            16'd2214: data <= 8'h00;
            16'd2215: data <= 8'hF8;
            16'd2216: data <= 8'h00;
            16'd2217: data <= 8'hF8;
            16'd2218: data <= 8'h00;
            16'd2219: data <= 8'hF8;
            16'd2220: data <= 8'h00;
            16'd2221: data <= 8'hF8;
            16'd2222: data <= 8'h00;
            16'd2223: data <= 8'hF8;
            16'd2224: data <= 8'h00;
            16'd2225: data <= 8'hF8;
            16'd2226: data <= 8'h00;
            16'd2227: data <= 8'hF8;
            16'd2228: data <= 8'h00;
            16'd2229: data <= 8'hF8;
            16'd2230: data <= 8'h00;
            16'd2231: data <= 8'hF8;
            16'd2232: data <= 8'h00;
            16'd2233: data <= 8'hF8;
            16'd2234: data <= 8'h00;
            16'd2235: data <= 8'hF8;
            16'd2236: data <= 8'h00;
            16'd2237: data <= 8'hF8;
            16'd2238: data <= 8'h00;
            16'd2239: data <= 8'hF8;
            16'd2240: data <= 8'hFF;
            16'd2241: data <= 8'hFF;
            16'd2242: data <= 8'h00;
            16'd2243: data <= 8'hF8;
            16'd2244: data <= 8'h00;
            16'd2245: data <= 8'hF8;
            16'd2246: data <= 8'h00;
            16'd2247: data <= 8'hF8;
            16'd2248: data <= 8'h00;
            16'd2249: data <= 8'hF8;
            16'd2250: data <= 8'h00;
            16'd2251: data <= 8'hF8;
            16'd2252: data <= 8'h00;
            16'd2253: data <= 8'hF8;
            16'd2254: data <= 8'h00;
            16'd2255: data <= 8'hF8;
            16'd2256: data <= 8'h00;
            16'd2257: data <= 8'hF8;
            16'd2258: data <= 8'h00;
            16'd2259: data <= 8'hF8;
            16'd2260: data <= 8'h00;
            16'd2261: data <= 8'hF8;
            16'd2262: data <= 8'h00;
            16'd2263: data <= 8'hF8;
            16'd2264: data <= 8'h00;
            16'd2265: data <= 8'hF8;
            16'd2266: data <= 8'h00;
            16'd2267: data <= 8'hF8;
            16'd2268: data <= 8'h00;
            16'd2269: data <= 8'hF8;
            16'd2270: data <= 8'h00;
            16'd2271: data <= 8'hF8;
            16'd2272: data <= 8'h00;
            16'd2273: data <= 8'hF8;
            16'd2274: data <= 8'h00;
            16'd2275: data <= 8'hF8;
            16'd2276: data <= 8'h00;
            16'd2277: data <= 8'hF8;
            16'd2278: data <= 8'h00;
            16'd2279: data <= 8'hF8;
            16'd2280: data <= 8'hFF;
            16'd2281: data <= 8'hFF;
            16'd2282: data <= 8'h00;
            16'd2283: data <= 8'hF8;
            16'd2284: data <= 8'h00;
            16'd2285: data <= 8'hF8;
            16'd2286: data <= 8'h00;
            16'd2287: data <= 8'hF8;
            16'd2288: data <= 8'h00;
            16'd2289: data <= 8'hF8;
            16'd2290: data <= 8'h00;
            16'd2291: data <= 8'hF8;
            16'd2292: data <= 8'h00;
            16'd2293: data <= 8'hF8;
            16'd2294: data <= 8'h00;
            16'd2295: data <= 8'hF8;
            16'd2296: data <= 8'h00;
            16'd2297: data <= 8'hF8;
            16'd2298: data <= 8'h00;
            16'd2299: data <= 8'hF8;
            16'd2300: data <= 8'h00;
            16'd2301: data <= 8'hF8;
            16'd2302: data <= 8'h00;
            16'd2303: data <= 8'hF8;
            16'd2304: data <= 8'h00;
            16'd2305: data <= 8'hF8;
            16'd2306: data <= 8'h00;
            16'd2307: data <= 8'hF8;
            16'd2308: data <= 8'h00;
            16'd2309: data <= 8'hF8;
            16'd2310: data <= 8'h00;
            16'd2311: data <= 8'hF8;
            16'd2312: data <= 8'h00;
            16'd2313: data <= 8'hF8;
            16'd2314: data <= 8'h00;
            16'd2315: data <= 8'hF8;
            16'd2316: data <= 8'h00;
            16'd2317: data <= 8'hF8;
            16'd2318: data <= 8'h00;
            16'd2319: data <= 8'hF8;
            16'd2320: data <= 8'hFF;
            16'd2321: data <= 8'hFF;
            16'd2322: data <= 8'h00;
            16'd2323: data <= 8'hF8;
            16'd2324: data <= 8'h00;
            16'd2325: data <= 8'hF8;
            16'd2326: data <= 8'h00;
            16'd2327: data <= 8'hF8;
            16'd2328: data <= 8'h00;
            16'd2329: data <= 8'hF8;
            16'd2330: data <= 8'h00;
            16'd2331: data <= 8'hF8;
            16'd2332: data <= 8'h00;
            16'd2333: data <= 8'hF8;
            16'd2334: data <= 8'h00;
            16'd2335: data <= 8'hF8;
            16'd2336: data <= 8'h00;
            16'd2337: data <= 8'hF8;
            16'd2338: data <= 8'h00;
            16'd2339: data <= 8'hF8;
            16'd2340: data <= 8'h00;
            16'd2341: data <= 8'hF8;
            16'd2342: data <= 8'h00;
            16'd2343: data <= 8'hF8;
            16'd2344: data <= 8'h00;
            16'd2345: data <= 8'hF8;
            16'd2346: data <= 8'h00;
            16'd2347: data <= 8'hF8;
            16'd2348: data <= 8'h00;
            16'd2349: data <= 8'hF8;
            16'd2350: data <= 8'h00;
            16'd2351: data <= 8'hF8;
            16'd2352: data <= 8'h00;
            16'd2353: data <= 8'hF8;
            16'd2354: data <= 8'h00;
            16'd2355: data <= 8'hF8;
            16'd2356: data <= 8'h00;
            16'd2357: data <= 8'hF8;
            16'd2358: data <= 8'h00;
            16'd2359: data <= 8'hF8;
            16'd2360: data <= 8'hFF;
            16'd2361: data <= 8'hFF;
            16'd2362: data <= 8'h00;
            16'd2363: data <= 8'hF8;
            16'd2364: data <= 8'h00;
            16'd2365: data <= 8'hF8;
            16'd2366: data <= 8'h00;
            16'd2367: data <= 8'hF8;
            16'd2368: data <= 8'h00;
            16'd2369: data <= 8'hF8;
            16'd2370: data <= 8'h00;
            16'd2371: data <= 8'hF8;
            16'd2372: data <= 8'h00;
            16'd2373: data <= 8'hF8;
            16'd2374: data <= 8'h00;
            16'd2375: data <= 8'hF8;
            16'd2376: data <= 8'h00;
            16'd2377: data <= 8'hF8;
            16'd2378: data <= 8'h00;
            16'd2379: data <= 8'hF8;
            16'd2380: data <= 8'h00;
            16'd2381: data <= 8'hF8;
            16'd2382: data <= 8'h00;
            16'd2383: data <= 8'hF8;
            16'd2384: data <= 8'h00;
            16'd2385: data <= 8'hF8;
            16'd2386: data <= 8'h00;
            16'd2387: data <= 8'hF8;
            16'd2388: data <= 8'h00;
            16'd2389: data <= 8'hF8;
            16'd2390: data <= 8'h00;
            16'd2391: data <= 8'hF8;
            16'd2392: data <= 8'h00;
            16'd2393: data <= 8'hF8;
            16'd2394: data <= 8'h00;
            16'd2395: data <= 8'hF8;
            16'd2396: data <= 8'h00;
            16'd2397: data <= 8'hF8;
            16'd2398: data <= 8'h00;
            16'd2399: data <= 8'hF8;
            16'd2400: data <= 8'hFF;
            16'd2401: data <= 8'hFF;
            16'd2402: data <= 8'h00;
            16'd2403: data <= 8'hF8;
            16'd2404: data <= 8'h00;
            16'd2405: data <= 8'hF8;
            16'd2406: data <= 8'h00;
            16'd2407: data <= 8'hF8;
            16'd2408: data <= 8'h00;
            16'd2409: data <= 8'hF8;
            16'd2410: data <= 8'h00;
            16'd2411: data <= 8'hF8;
            16'd2412: data <= 8'h00;
            16'd2413: data <= 8'hF8;
            16'd2414: data <= 8'h00;
            16'd2415: data <= 8'hF8;
            16'd2416: data <= 8'h00;
            16'd2417: data <= 8'hF8;
            16'd2418: data <= 8'h00;
            16'd2419: data <= 8'hF8;
            16'd2420: data <= 8'h00;
            16'd2421: data <= 8'hF8;
            16'd2422: data <= 8'h00;
            16'd2423: data <= 8'hF8;
            16'd2424: data <= 8'h00;
            16'd2425: data <= 8'hF8;
            16'd2426: data <= 8'h00;
            16'd2427: data <= 8'hF8;
            16'd2428: data <= 8'h00;
            16'd2429: data <= 8'hF8;
            16'd2430: data <= 8'h00;
            16'd2431: data <= 8'hF8;
            16'd2432: data <= 8'h00;
            16'd2433: data <= 8'hF8;
            16'd2434: data <= 8'h00;
            16'd2435: data <= 8'hF8;
            16'd2436: data <= 8'h00;
            16'd2437: data <= 8'hF8;
            16'd2438: data <= 8'h00;
            16'd2439: data <= 8'hF8;
            16'd2440: data <= 8'hFF;
            16'd2441: data <= 8'hFF;
            16'd2442: data <= 8'h00;
            16'd2443: data <= 8'hF8;
            16'd2444: data <= 8'h00;
            16'd2445: data <= 8'hF8;
            16'd2446: data <= 8'h00;
            16'd2447: data <= 8'hF8;
            16'd2448: data <= 8'h00;
            16'd2449: data <= 8'hF8;
            16'd2450: data <= 8'h00;
            16'd2451: data <= 8'hF8;
            16'd2452: data <= 8'h00;
            16'd2453: data <= 8'hF8;
            16'd2454: data <= 8'h00;
            16'd2455: data <= 8'hF8;
            16'd2456: data <= 8'h00;
            16'd2457: data <= 8'hF8;
            16'd2458: data <= 8'h00;
            16'd2459: data <= 8'hF8;
            16'd2460: data <= 8'h00;
            16'd2461: data <= 8'hF8;
            16'd2462: data <= 8'h00;
            16'd2463: data <= 8'hF8;
            16'd2464: data <= 8'h00;
            16'd2465: data <= 8'hF8;
            16'd2466: data <= 8'h00;
            16'd2467: data <= 8'hF8;
            16'd2468: data <= 8'h00;
            16'd2469: data <= 8'hF8;
            16'd2470: data <= 8'h00;
            16'd2471: data <= 8'hF8;
            16'd2472: data <= 8'h00;
            16'd2473: data <= 8'hF8;
            16'd2474: data <= 8'h00;
            16'd2475: data <= 8'hF8;
            16'd2476: data <= 8'h00;
            16'd2477: data <= 8'hF8;
            16'd2478: data <= 8'h00;
            16'd2479: data <= 8'hF8;
            16'd2480: data <= 8'hFF;
            16'd2481: data <= 8'hFF;
            16'd2482: data <= 8'h00;
            16'd2483: data <= 8'hF8;
            16'd2484: data <= 8'h00;
            16'd2485: data <= 8'hF8;
            16'd2486: data <= 8'h00;
            16'd2487: data <= 8'hF8;
            16'd2488: data <= 8'h00;
            16'd2489: data <= 8'hF8;
            16'd2490: data <= 8'h00;
            16'd2491: data <= 8'hF8;
            16'd2492: data <= 8'h00;
            16'd2493: data <= 8'hF8;
            16'd2494: data <= 8'h00;
            16'd2495: data <= 8'hF8;
            16'd2496: data <= 8'h00;
            16'd2497: data <= 8'hF8;
            16'd2498: data <= 8'h00;
            16'd2499: data <= 8'hF8;
            16'd2500: data <= 8'h00;
            16'd2501: data <= 8'hF8;
            16'd2502: data <= 8'h00;
            16'd2503: data <= 8'hF8;
            16'd2504: data <= 8'h00;
            16'd2505: data <= 8'hF8;
            16'd2506: data <= 8'h00;
            16'd2507: data <= 8'hF8;
            16'd2508: data <= 8'h00;
            16'd2509: data <= 8'hF8;
            16'd2510: data <= 8'h00;
            16'd2511: data <= 8'hF8;
            16'd2512: data <= 8'h00;
            16'd2513: data <= 8'hF8;
            16'd2514: data <= 8'h00;
            16'd2515: data <= 8'hF8;
            16'd2516: data <= 8'h00;
            16'd2517: data <= 8'hF8;
            16'd2518: data <= 8'h00;
            16'd2519: data <= 8'hF8;
            16'd2520: data <= 8'hFF;
            16'd2521: data <= 8'hFF;
            16'd2522: data <= 8'h00;
            16'd2523: data <= 8'hF8;
            16'd2524: data <= 8'h00;
            16'd2525: data <= 8'hF8;
            16'd2526: data <= 8'h00;
            16'd2527: data <= 8'hF8;
            16'd2528: data <= 8'h00;
            16'd2529: data <= 8'hF8;
            16'd2530: data <= 8'h00;
            16'd2531: data <= 8'hF8;
            16'd2532: data <= 8'h00;
            16'd2533: data <= 8'hF8;
            16'd2534: data <= 8'h00;
            16'd2535: data <= 8'hF8;
            16'd2536: data <= 8'h00;
            16'd2537: data <= 8'hF8;
            16'd2538: data <= 8'h00;
            16'd2539: data <= 8'hF8;
            16'd2540: data <= 8'h00;
            16'd2541: data <= 8'hF8;
            16'd2542: data <= 8'h00;
            16'd2543: data <= 8'hF8;
            16'd2544: data <= 8'h00;
            16'd2545: data <= 8'hF8;
            16'd2546: data <= 8'h00;
            16'd2547: data <= 8'hF8;
            16'd2548: data <= 8'h00;
            16'd2549: data <= 8'hF8;
            16'd2550: data <= 8'h00;
            16'd2551: data <= 8'hF8;
            16'd2552: data <= 8'h00;
            16'd2553: data <= 8'hF8;
            16'd2554: data <= 8'h00;
            16'd2555: data <= 8'hF8;
            16'd2556: data <= 8'h00;
            16'd2557: data <= 8'hF8;
            16'd2558: data <= 8'h00;
            16'd2559: data <= 8'hF8;
            16'd2560: data <= 8'hFF;
            16'd2561: data <= 8'hFF;
            16'd2562: data <= 8'h00;
            16'd2563: data <= 8'hF8;
            16'd2564: data <= 8'h00;
            16'd2565: data <= 8'hF8;
            16'd2566: data <= 8'h00;
            16'd2567: data <= 8'hF8;
            16'd2568: data <= 8'h00;
            16'd2569: data <= 8'hF8;
            16'd2570: data <= 8'h00;
            16'd2571: data <= 8'hF8;
            16'd2572: data <= 8'h00;
            16'd2573: data <= 8'hF8;
            16'd2574: data <= 8'h00;
            16'd2575: data <= 8'hF8;
            16'd2576: data <= 8'h00;
            16'd2577: data <= 8'hF8;
            16'd2578: data <= 8'h00;
            16'd2579: data <= 8'hF8;
            16'd2580: data <= 8'h00;
            16'd2581: data <= 8'hF8;
            16'd2582: data <= 8'h00;
            16'd2583: data <= 8'hF8;
            16'd2584: data <= 8'h00;
            16'd2585: data <= 8'hF8;
            16'd2586: data <= 8'h00;
            16'd2587: data <= 8'hF8;
            16'd2588: data <= 8'h00;
            16'd2589: data <= 8'hF8;
            16'd2590: data <= 8'h00;
            16'd2591: data <= 8'hF8;
            16'd2592: data <= 8'h00;
            16'd2593: data <= 8'hF8;
            16'd2594: data <= 8'h00;
            16'd2595: data <= 8'hF8;
            16'd2596: data <= 8'h00;
            16'd2597: data <= 8'hF8;
            16'd2598: data <= 8'h00;
            16'd2599: data <= 8'hF8;
            16'd2600: data <= 8'hFF;
            16'd2601: data <= 8'hFF;
            16'd2602: data <= 8'h00;
            16'd2603: data <= 8'hF8;
            16'd2604: data <= 8'h00;
            16'd2605: data <= 8'hF8;
            16'd2606: data <= 8'h00;
            16'd2607: data <= 8'hF8;
            16'd2608: data <= 8'h00;
            16'd2609: data <= 8'hF8;
            16'd2610: data <= 8'h00;
            16'd2611: data <= 8'hF8;
            16'd2612: data <= 8'h00;
            16'd2613: data <= 8'hF8;
            16'd2614: data <= 8'h00;
            16'd2615: data <= 8'hF8;
            16'd2616: data <= 8'h00;
            16'd2617: data <= 8'hF8;
            16'd2618: data <= 8'h00;
            16'd2619: data <= 8'hF8;
            16'd2620: data <= 8'h00;
            16'd2621: data <= 8'hF8;
            16'd2622: data <= 8'h00;
            16'd2623: data <= 8'hF8;
            16'd2624: data <= 8'h00;
            16'd2625: data <= 8'hF8;
            16'd2626: data <= 8'h00;
            16'd2627: data <= 8'hF8;
            16'd2628: data <= 8'h00;
            16'd2629: data <= 8'hF8;
            16'd2630: data <= 8'h00;
            16'd2631: data <= 8'hF8;
            16'd2632: data <= 8'h00;
            16'd2633: data <= 8'hF8;
            16'd2634: data <= 8'h00;
            16'd2635: data <= 8'hF8;
            16'd2636: data <= 8'h00;
            16'd2637: data <= 8'hF8;
            16'd2638: data <= 8'h00;
            16'd2639: data <= 8'hF8;
            16'd2640: data <= 8'hFF;
            16'd2641: data <= 8'hFF;
            16'd2642: data <= 8'h00;
            16'd2643: data <= 8'hF8;
            16'd2644: data <= 8'h00;
            16'd2645: data <= 8'hF8;
            16'd2646: data <= 8'h00;
            16'd2647: data <= 8'hF8;
            16'd2648: data <= 8'h00;
            16'd2649: data <= 8'hF8;
            16'd2650: data <= 8'h00;
            16'd2651: data <= 8'hF8;
            16'd2652: data <= 8'h00;
            16'd2653: data <= 8'hF8;
            16'd2654: data <= 8'h00;
            16'd2655: data <= 8'hF8;
            16'd2656: data <= 8'h00;
            16'd2657: data <= 8'hF8;
            16'd2658: data <= 8'h00;
            16'd2659: data <= 8'hF8;
            16'd2660: data <= 8'h00;
            16'd2661: data <= 8'hF8;
            16'd2662: data <= 8'h00;
            16'd2663: data <= 8'hF8;
            16'd2664: data <= 8'h00;
            16'd2665: data <= 8'hF8;
            16'd2666: data <= 8'h00;
            16'd2667: data <= 8'hF8;
            16'd2668: data <= 8'h00;
            16'd2669: data <= 8'hF8;
            16'd2670: data <= 8'h00;
            16'd2671: data <= 8'hF8;
            16'd2672: data <= 8'h00;
            16'd2673: data <= 8'hF8;
            16'd2674: data <= 8'h00;
            16'd2675: data <= 8'hF8;
            16'd2676: data <= 8'h00;
            16'd2677: data <= 8'hF8;
            16'd2678: data <= 8'h00;
            16'd2679: data <= 8'hF8;
            16'd2680: data <= 8'hFF;
            16'd2681: data <= 8'hFF;
            16'd2682: data <= 8'h00;
            16'd2683: data <= 8'hF8;
            16'd2684: data <= 8'h00;
            16'd2685: data <= 8'hF8;
            16'd2686: data <= 8'h00;
            16'd2687: data <= 8'hF8;
            16'd2688: data <= 8'h00;
            16'd2689: data <= 8'hF8;
            16'd2690: data <= 8'h00;
            16'd2691: data <= 8'hF8;
            16'd2692: data <= 8'h00;
            16'd2693: data <= 8'hF8;
            16'd2694: data <= 8'h00;
            16'd2695: data <= 8'hF8;
            16'd2696: data <= 8'h00;
            16'd2697: data <= 8'hF8;
            16'd2698: data <= 8'h00;
            16'd2699: data <= 8'hF8;
            16'd2700: data <= 8'h00;
            16'd2701: data <= 8'hF8;
            16'd2702: data <= 8'h00;
            16'd2703: data <= 8'hF8;
            16'd2704: data <= 8'h00;
            16'd2705: data <= 8'hF8;
            16'd2706: data <= 8'h00;
            16'd2707: data <= 8'hF8;
            16'd2708: data <= 8'h00;
            16'd2709: data <= 8'hF8;
            16'd2710: data <= 8'h00;
            16'd2711: data <= 8'hF8;
            16'd2712: data <= 8'h00;
            16'd2713: data <= 8'hF8;
            16'd2714: data <= 8'h00;
            16'd2715: data <= 8'hF8;
            16'd2716: data <= 8'h00;
            16'd2717: data <= 8'hF8;
            16'd2718: data <= 8'h00;
            16'd2719: data <= 8'hF8;
            16'd2720: data <= 8'hFF;
            16'd2721: data <= 8'hFF;
            16'd2722: data <= 8'h00;
            16'd2723: data <= 8'hF8;
            16'd2724: data <= 8'h00;
            16'd2725: data <= 8'hF8;
            16'd2726: data <= 8'h00;
            16'd2727: data <= 8'hF8;
            16'd2728: data <= 8'h00;
            16'd2729: data <= 8'hF8;
            16'd2730: data <= 8'h00;
            16'd2731: data <= 8'hF8;
            16'd2732: data <= 8'h00;
            16'd2733: data <= 8'hF8;
            16'd2734: data <= 8'h00;
            16'd2735: data <= 8'hF8;
            16'd2736: data <= 8'h00;
            16'd2737: data <= 8'hF8;
            16'd2738: data <= 8'h00;
            16'd2739: data <= 8'hF8;
            16'd2740: data <= 8'h00;
            16'd2741: data <= 8'hF8;
            16'd2742: data <= 8'h00;
            16'd2743: data <= 8'hF8;
            16'd2744: data <= 8'h00;
            16'd2745: data <= 8'hF8;
            16'd2746: data <= 8'h00;
            16'd2747: data <= 8'hF8;
            16'd2748: data <= 8'h00;
            16'd2749: data <= 8'hF8;
            16'd2750: data <= 8'h00;
            16'd2751: data <= 8'hF8;
            16'd2752: data <= 8'h00;
            16'd2753: data <= 8'hF8;
            16'd2754: data <= 8'h00;
            16'd2755: data <= 8'hF8;
            16'd2756: data <= 8'h00;
            16'd2757: data <= 8'hF8;
            16'd2758: data <= 8'h00;
            16'd2759: data <= 8'hF8;
            16'd2760: data <= 8'hFF;
            16'd2761: data <= 8'hFF;
            16'd2762: data <= 8'h00;
            16'd2763: data <= 8'hF8;
            16'd2764: data <= 8'h00;
            16'd2765: data <= 8'hF8;
            16'd2766: data <= 8'h00;
            16'd2767: data <= 8'hF8;
            16'd2768: data <= 8'h00;
            16'd2769: data <= 8'hF8;
            16'd2770: data <= 8'h00;
            16'd2771: data <= 8'hF8;
            16'd2772: data <= 8'h00;
            16'd2773: data <= 8'hF8;
            16'd2774: data <= 8'h00;
            16'd2775: data <= 8'hF8;
            16'd2776: data <= 8'h00;
            16'd2777: data <= 8'hF8;
            16'd2778: data <= 8'h00;
            16'd2779: data <= 8'hF8;
            16'd2780: data <= 8'h00;
            16'd2781: data <= 8'hF8;
            16'd2782: data <= 8'h00;
            16'd2783: data <= 8'hF8;
            16'd2784: data <= 8'h00;
            16'd2785: data <= 8'hF8;
            16'd2786: data <= 8'h00;
            16'd2787: data <= 8'hF8;
            16'd2788: data <= 8'h00;
            16'd2789: data <= 8'hF8;
            16'd2790: data <= 8'h00;
            16'd2791: data <= 8'hF8;
            16'd2792: data <= 8'h00;
            16'd2793: data <= 8'hF8;
            16'd2794: data <= 8'h00;
            16'd2795: data <= 8'hF8;
            16'd2796: data <= 8'h00;
            16'd2797: data <= 8'hF8;
            16'd2798: data <= 8'h00;
            16'd2799: data <= 8'hF8;
            16'd2800: data <= 8'hFF;
            16'd2801: data <= 8'hFF;
            16'd2802: data <= 8'h00;
            16'd2803: data <= 8'hF8;
            16'd2804: data <= 8'h00;
            16'd2805: data <= 8'hF8;
            16'd2806: data <= 8'h00;
            16'd2807: data <= 8'hF8;
            16'd2808: data <= 8'h00;
            16'd2809: data <= 8'hF8;
            16'd2810: data <= 8'h00;
            16'd2811: data <= 8'hF8;
            16'd2812: data <= 8'h00;
            16'd2813: data <= 8'hF8;
            16'd2814: data <= 8'h00;
            16'd2815: data <= 8'hF8;
            16'd2816: data <= 8'h00;
            16'd2817: data <= 8'hF8;
            16'd2818: data <= 8'h00;
            16'd2819: data <= 8'hF8;
            16'd2820: data <= 8'h00;
            16'd2821: data <= 8'hF8;
            16'd2822: data <= 8'h00;
            16'd2823: data <= 8'hF8;
            16'd2824: data <= 8'h00;
            16'd2825: data <= 8'hF8;
            16'd2826: data <= 8'h00;
            16'd2827: data <= 8'hF8;
            16'd2828: data <= 8'h00;
            16'd2829: data <= 8'hF8;
            16'd2830: data <= 8'h00;
            16'd2831: data <= 8'hF8;
            16'd2832: data <= 8'h00;
            16'd2833: data <= 8'hF8;
            16'd2834: data <= 8'h00;
            16'd2835: data <= 8'hF8;
            16'd2836: data <= 8'h00;
            16'd2837: data <= 8'hF8;
            16'd2838: data <= 8'h00;
            16'd2839: data <= 8'hF8;
            16'd2840: data <= 8'hFF;
            16'd2841: data <= 8'hFF;
            16'd2842: data <= 8'h00;
            16'd2843: data <= 8'hF8;
            16'd2844: data <= 8'h00;
            16'd2845: data <= 8'hF8;
            16'd2846: data <= 8'h00;
            16'd2847: data <= 8'hF8;
            16'd2848: data <= 8'h00;
            16'd2849: data <= 8'hF8;
            16'd2850: data <= 8'h00;
            16'd2851: data <= 8'hF8;
            16'd2852: data <= 8'h00;
            16'd2853: data <= 8'hF8;
            16'd2854: data <= 8'h00;
            16'd2855: data <= 8'hF8;
            16'd2856: data <= 8'h00;
            16'd2857: data <= 8'hF8;
            16'd2858: data <= 8'h00;
            16'd2859: data <= 8'hF8;
            16'd2860: data <= 8'h00;
            16'd2861: data <= 8'hF8;
            16'd2862: data <= 8'h00;
            16'd2863: data <= 8'hF8;
            16'd2864: data <= 8'h00;
            16'd2865: data <= 8'hF8;
            16'd2866: data <= 8'h00;
            16'd2867: data <= 8'hF8;
            16'd2868: data <= 8'h00;
            16'd2869: data <= 8'hF8;
            16'd2870: data <= 8'h00;
            16'd2871: data <= 8'hF8;
            16'd2872: data <= 8'h00;
            16'd2873: data <= 8'hF8;
            16'd2874: data <= 8'h00;
            16'd2875: data <= 8'hF8;
            16'd2876: data <= 8'h00;
            16'd2877: data <= 8'hF8;
            16'd2878: data <= 8'h00;
            16'd2879: data <= 8'hF8;
            16'd2880: data <= 8'hFF;
            16'd2881: data <= 8'hFF;
            16'd2882: data <= 8'h00;
            16'd2883: data <= 8'hF8;
            16'd2884: data <= 8'h00;
            16'd2885: data <= 8'hF8;
            16'd2886: data <= 8'h00;
            16'd2887: data <= 8'hF8;
            16'd2888: data <= 8'h00;
            16'd2889: data <= 8'hF8;
            16'd2890: data <= 8'h00;
            16'd2891: data <= 8'hF8;
            16'd2892: data <= 8'h00;
            16'd2893: data <= 8'hF8;
            16'd2894: data <= 8'h00;
            16'd2895: data <= 8'hF8;
            16'd2896: data <= 8'h00;
            16'd2897: data <= 8'hF8;
            16'd2898: data <= 8'h00;
            16'd2899: data <= 8'hF8;
            16'd2900: data <= 8'h00;
            16'd2901: data <= 8'hF8;
            16'd2902: data <= 8'h00;
            16'd2903: data <= 8'hF8;
            16'd2904: data <= 8'h00;
            16'd2905: data <= 8'hF8;
            16'd2906: data <= 8'h00;
            16'd2907: data <= 8'hF8;
            16'd2908: data <= 8'h00;
            16'd2909: data <= 8'hF8;
            16'd2910: data <= 8'h00;
            16'd2911: data <= 8'hF8;
            16'd2912: data <= 8'h00;
            16'd2913: data <= 8'hF8;
            16'd2914: data <= 8'h00;
            16'd2915: data <= 8'hF8;
            16'd2916: data <= 8'h00;
            16'd2917: data <= 8'hF8;
            16'd2918: data <= 8'h00;
            16'd2919: data <= 8'hF8;
            16'd2920: data <= 8'hFF;
            16'd2921: data <= 8'hFF;
            16'd2922: data <= 8'h00;
            16'd2923: data <= 8'hF8;
            16'd2924: data <= 8'h00;
            16'd2925: data <= 8'hF8;
            16'd2926: data <= 8'h00;
            16'd2927: data <= 8'hF8;
            16'd2928: data <= 8'h00;
            16'd2929: data <= 8'hF8;
            16'd2930: data <= 8'h00;
            16'd2931: data <= 8'hF8;
            16'd2932: data <= 8'h00;
            16'd2933: data <= 8'hF8;
            16'd2934: data <= 8'h00;
            16'd2935: data <= 8'hF8;
            16'd2936: data <= 8'h00;
            16'd2937: data <= 8'hF8;
            16'd2938: data <= 8'h00;
            16'd2939: data <= 8'hF8;
            16'd2940: data <= 8'h00;
            16'd2941: data <= 8'hF8;
            16'd2942: data <= 8'h00;
            16'd2943: data <= 8'hF8;
            16'd2944: data <= 8'h00;
            16'd2945: data <= 8'hF8;
            16'd2946: data <= 8'h00;
            16'd2947: data <= 8'hF8;
            16'd2948: data <= 8'h00;
            16'd2949: data <= 8'hF8;
            16'd2950: data <= 8'h00;
            16'd2951: data <= 8'hF8;
            16'd2952: data <= 8'h00;
            16'd2953: data <= 8'hF8;
            16'd2954: data <= 8'h00;
            16'd2955: data <= 8'hF8;
            16'd2956: data <= 8'h00;
            16'd2957: data <= 8'hF8;
            16'd2958: data <= 8'h00;
            16'd2959: data <= 8'hF8;
            16'd2960: data <= 8'hFF;
            16'd2961: data <= 8'hFF;
            16'd2962: data <= 8'h00;
            16'd2963: data <= 8'hF8;
            16'd2964: data <= 8'h00;
            16'd2965: data <= 8'hF8;
            16'd2966: data <= 8'h00;
            16'd2967: data <= 8'hF8;
            16'd2968: data <= 8'h00;
            16'd2969: data <= 8'hF8;
            16'd2970: data <= 8'h00;
            16'd2971: data <= 8'hF8;
            16'd2972: data <= 8'h00;
            16'd2973: data <= 8'hF8;
            16'd2974: data <= 8'h00;
            16'd2975: data <= 8'hF8;
            16'd2976: data <= 8'h00;
            16'd2977: data <= 8'hF8;
            16'd2978: data <= 8'h00;
            16'd2979: data <= 8'hF8;
            16'd2980: data <= 8'h00;
            16'd2981: data <= 8'hF8;
            16'd2982: data <= 8'h00;
            16'd2983: data <= 8'hF8;
            16'd2984: data <= 8'h00;
            16'd2985: data <= 8'hF8;
            16'd2986: data <= 8'h00;
            16'd2987: data <= 8'hF8;
            16'd2988: data <= 8'h00;
            16'd2989: data <= 8'hF8;
            16'd2990: data <= 8'h00;
            16'd2991: data <= 8'hF8;
            16'd2992: data <= 8'h00;
            16'd2993: data <= 8'hF8;
            16'd2994: data <= 8'h00;
            16'd2995: data <= 8'hF8;
            16'd2996: data <= 8'h00;
            16'd2997: data <= 8'hF8;
            16'd2998: data <= 8'h00;
            16'd2999: data <= 8'hF8;
            16'd3000: data <= 8'hFF;
            16'd3001: data <= 8'hFF;
            16'd3002: data <= 8'h00;
            16'd3003: data <= 8'hF8;
            16'd3004: data <= 8'h00;
            16'd3005: data <= 8'hF8;
            16'd3006: data <= 8'h00;
            16'd3007: data <= 8'hF8;
            16'd3008: data <= 8'h00;
            16'd3009: data <= 8'hF8;
            16'd3010: data <= 8'h00;
            16'd3011: data <= 8'hF8;
            16'd3012: data <= 8'h00;
            16'd3013: data <= 8'hF8;
            16'd3014: data <= 8'h00;
            16'd3015: data <= 8'hF8;
            16'd3016: data <= 8'h00;
            16'd3017: data <= 8'hF8;
            16'd3018: data <= 8'h00;
            16'd3019: data <= 8'hF8;
            16'd3020: data <= 8'h00;
            16'd3021: data <= 8'hF8;
            16'd3022: data <= 8'h00;
            16'd3023: data <= 8'hF8;
            16'd3024: data <= 8'h00;
            16'd3025: data <= 8'hF8;
            16'd3026: data <= 8'h00;
            16'd3027: data <= 8'hF8;
            16'd3028: data <= 8'h00;
            16'd3029: data <= 8'hF8;
            16'd3030: data <= 8'h00;
            16'd3031: data <= 8'hF8;
            16'd3032: data <= 8'h00;
            16'd3033: data <= 8'hF8;
            16'd3034: data <= 8'h00;
            16'd3035: data <= 8'hF8;
            16'd3036: data <= 8'h00;
            16'd3037: data <= 8'hF8;
            16'd3038: data <= 8'h00;
            16'd3039: data <= 8'hF8;
            16'd3040: data <= 8'hFF;
            16'd3041: data <= 8'hFF;
            16'd3042: data <= 8'h00;
            16'd3043: data <= 8'hF8;
            16'd3044: data <= 8'h00;
            16'd3045: data <= 8'hF8;
            16'd3046: data <= 8'h00;
            16'd3047: data <= 8'hF8;
            16'd3048: data <= 8'h00;
            16'd3049: data <= 8'hF8;
            16'd3050: data <= 8'h00;
            16'd3051: data <= 8'hF8;
            16'd3052: data <= 8'h00;
            16'd3053: data <= 8'hF8;
            16'd3054: data <= 8'h00;
            16'd3055: data <= 8'hF8;
            16'd3056: data <= 8'h00;
            16'd3057: data <= 8'hF8;
            16'd3058: data <= 8'h00;
            16'd3059: data <= 8'hF8;
            16'd3060: data <= 8'h00;
            16'd3061: data <= 8'hF8;
            16'd3062: data <= 8'h00;
            16'd3063: data <= 8'hF8;
            16'd3064: data <= 8'h00;
            16'd3065: data <= 8'hF8;
            16'd3066: data <= 8'h00;
            16'd3067: data <= 8'hF8;
            16'd3068: data <= 8'h00;
            16'd3069: data <= 8'hF8;
            16'd3070: data <= 8'h00;
            16'd3071: data <= 8'hF8;
            16'd3072: data <= 8'h00;
            16'd3073: data <= 8'hF8;
            16'd3074: data <= 8'h00;
            16'd3075: data <= 8'hF8;
            16'd3076: data <= 8'h00;
            16'd3077: data <= 8'hF8;
            16'd3078: data <= 8'h00;
            16'd3079: data <= 8'hF8;
            16'd3080: data <= 8'hFF;
            16'd3081: data <= 8'hFF;
            16'd3082: data <= 8'h00;
            16'd3083: data <= 8'hF8;
            16'd3084: data <= 8'h00;
            16'd3085: data <= 8'hF8;
            16'd3086: data <= 8'h00;
            16'd3087: data <= 8'hF8;
            16'd3088: data <= 8'h00;
            16'd3089: data <= 8'hF8;
            16'd3090: data <= 8'h00;
            16'd3091: data <= 8'hF8;
            16'd3092: data <= 8'h00;
            16'd3093: data <= 8'hF8;
            16'd3094: data <= 8'h00;
            16'd3095: data <= 8'hF8;
            16'd3096: data <= 8'h00;
            16'd3097: data <= 8'hF8;
            16'd3098: data <= 8'h00;
            16'd3099: data <= 8'hF8;
            16'd3100: data <= 8'h00;
            16'd3101: data <= 8'hF8;
            16'd3102: data <= 8'h00;
            16'd3103: data <= 8'hF8;
            16'd3104: data <= 8'h00;
            16'd3105: data <= 8'hF8;
            16'd3106: data <= 8'h00;
            16'd3107: data <= 8'hF8;
            16'd3108: data <= 8'h00;
            16'd3109: data <= 8'hF8;
            16'd3110: data <= 8'h00;
            16'd3111: data <= 8'hF8;
            16'd3112: data <= 8'h00;
            16'd3113: data <= 8'hF8;
            16'd3114: data <= 8'h00;
            16'd3115: data <= 8'hF8;
            16'd3116: data <= 8'h00;
            16'd3117: data <= 8'hF8;
            16'd3118: data <= 8'h00;
            16'd3119: data <= 8'hF8;
            16'd3120: data <= 8'hFF;
            16'd3121: data <= 8'hFF;
            16'd3122: data <= 8'h00;
            16'd3123: data <= 8'hF8;
            16'd3124: data <= 8'h00;
            16'd3125: data <= 8'hF8;
            16'd3126: data <= 8'h00;
            16'd3127: data <= 8'hF8;
            16'd3128: data <= 8'h00;
            16'd3129: data <= 8'hF8;
            16'd3130: data <= 8'h00;
            16'd3131: data <= 8'hF8;
            16'd3132: data <= 8'h00;
            16'd3133: data <= 8'hF8;
            16'd3134: data <= 8'h00;
            16'd3135: data <= 8'hF8;
            16'd3136: data <= 8'h00;
            16'd3137: data <= 8'hF8;
            16'd3138: data <= 8'h00;
            16'd3139: data <= 8'hF8;
            16'd3140: data <= 8'h00;
            16'd3141: data <= 8'hF8;
            16'd3142: data <= 8'h00;
            16'd3143: data <= 8'hF8;
            16'd3144: data <= 8'h00;
            16'd3145: data <= 8'hF8;
            16'd3146: data <= 8'h00;
            16'd3147: data <= 8'hF8;
            16'd3148: data <= 8'h00;
            16'd3149: data <= 8'hF8;
            16'd3150: data <= 8'h00;
            16'd3151: data <= 8'hF8;
            16'd3152: data <= 8'h00;
            16'd3153: data <= 8'hF8;
            16'd3154: data <= 8'h00;
            16'd3155: data <= 8'hF8;
            16'd3156: data <= 8'h00;
            16'd3157: data <= 8'hF8;
            16'd3158: data <= 8'h00;
            16'd3159: data <= 8'hF8;
            16'd3160: data <= 8'hFF;
            16'd3161: data <= 8'hFF;
            16'd3162: data <= 8'h00;
            16'd3163: data <= 8'hF8;
            16'd3164: data <= 8'h00;
            16'd3165: data <= 8'hF8;
            16'd3166: data <= 8'h00;
            16'd3167: data <= 8'hF8;
            16'd3168: data <= 8'h00;
            16'd3169: data <= 8'hF8;
            16'd3170: data <= 8'h00;
            16'd3171: data <= 8'hF8;
            16'd3172: data <= 8'h00;
            16'd3173: data <= 8'hF8;
            16'd3174: data <= 8'h00;
            16'd3175: data <= 8'hF8;
            16'd3176: data <= 8'h00;
            16'd3177: data <= 8'hF8;
            16'd3178: data <= 8'h00;
            16'd3179: data <= 8'hF8;
            16'd3180: data <= 8'h00;
            16'd3181: data <= 8'hF8;
            16'd3182: data <= 8'h00;
            16'd3183: data <= 8'hF8;
            16'd3184: data <= 8'h00;
            16'd3185: data <= 8'hF8;
            16'd3186: data <= 8'h00;
            16'd3187: data <= 8'hF8;
            16'd3188: data <= 8'h00;
            16'd3189: data <= 8'hF8;
            16'd3190: data <= 8'h00;
            16'd3191: data <= 8'hF8;
            16'd3192: data <= 8'h00;
            16'd3193: data <= 8'hF8;
            16'd3194: data <= 8'h00;
            16'd3195: data <= 8'hF8;
            16'd3196: data <= 8'h00;
            16'd3197: data <= 8'hF8;
            16'd3198: data <= 8'h00;
            16'd3199: data <= 8'hF8;
            16'd3200: data <= 8'hFF;
            16'd3201: data <= 8'hFF;
            16'd3202: data <= 8'h00;
            16'd3203: data <= 8'hF8;
            16'd3204: data <= 8'h00;
            16'd3205: data <= 8'hF8;
            16'd3206: data <= 8'h00;
            16'd3207: data <= 8'hF8;
            16'd3208: data <= 8'h00;
            16'd3209: data <= 8'hF8;
            16'd3210: data <= 8'h00;
            16'd3211: data <= 8'hF8;
            16'd3212: data <= 8'h00;
            16'd3213: data <= 8'hF8;
            16'd3214: data <= 8'h00;
            16'd3215: data <= 8'hF8;
            16'd3216: data <= 8'h00;
            16'd3217: data <= 8'hF8;
            16'd3218: data <= 8'h00;
            16'd3219: data <= 8'hF8;
            16'd3220: data <= 8'h00;
            16'd3221: data <= 8'hF8;
            16'd3222: data <= 8'h00;
            16'd3223: data <= 8'hF8;
            16'd3224: data <= 8'h00;
            16'd3225: data <= 8'hF8;
            16'd3226: data <= 8'h00;
            16'd3227: data <= 8'hF8;
            16'd3228: data <= 8'h00;
            16'd3229: data <= 8'hF8;
            16'd3230: data <= 8'h00;
            16'd3231: data <= 8'hF8;
            16'd3232: data <= 8'h00;
            16'd3233: data <= 8'hF8;
            16'd3234: data <= 8'h00;
            16'd3235: data <= 8'hF8;
            16'd3236: data <= 8'h00;
            16'd3237: data <= 8'hF8;
            16'd3238: data <= 8'h00;
            16'd3239: data <= 8'hF8;
            16'd3240: data <= 8'hFF;
            16'd3241: data <= 8'hFF;
            16'd3242: data <= 8'h00;
            16'd3243: data <= 8'hF8;
            16'd3244: data <= 8'h00;
            16'd3245: data <= 8'hF8;
            16'd3246: data <= 8'h00;
            16'd3247: data <= 8'hF8;
            16'd3248: data <= 8'h00;
            16'd3249: data <= 8'hF8;
            16'd3250: data <= 8'h00;
            16'd3251: data <= 8'hF8;
            16'd3252: data <= 8'h00;
            16'd3253: data <= 8'hF8;
            16'd3254: data <= 8'h00;
            16'd3255: data <= 8'hF8;
            16'd3256: data <= 8'h00;
            16'd3257: data <= 8'hF8;
            16'd3258: data <= 8'h00;
            16'd3259: data <= 8'hF8;
            16'd3260: data <= 8'h00;
            16'd3261: data <= 8'hF8;
            16'd3262: data <= 8'h00;
            16'd3263: data <= 8'hF8;
            16'd3264: data <= 8'h00;
            16'd3265: data <= 8'hF8;
            16'd3266: data <= 8'h00;
            16'd3267: data <= 8'hF8;
            16'd3268: data <= 8'h00;
            16'd3269: data <= 8'hF8;
            16'd3270: data <= 8'h00;
            16'd3271: data <= 8'hF8;
            16'd3272: data <= 8'h00;
            16'd3273: data <= 8'hF8;
            16'd3274: data <= 8'h00;
            16'd3275: data <= 8'hF8;
            16'd3276: data <= 8'h00;
            16'd3277: data <= 8'hF8;
            16'd3278: data <= 8'h00;
            16'd3279: data <= 8'hF8;
            16'd3280: data <= 8'hFF;
            16'd3281: data <= 8'hFF;
            16'd3282: data <= 8'h00;
            16'd3283: data <= 8'hF8;
            16'd3284: data <= 8'h00;
            16'd3285: data <= 8'hF8;
            16'd3286: data <= 8'h00;
            16'd3287: data <= 8'hF8;
            16'd3288: data <= 8'h00;
            16'd3289: data <= 8'hF8;
            16'd3290: data <= 8'h00;
            16'd3291: data <= 8'hF8;
            16'd3292: data <= 8'h00;
            16'd3293: data <= 8'hF8;
            16'd3294: data <= 8'h00;
            16'd3295: data <= 8'hF8;
            16'd3296: data <= 8'h00;
            16'd3297: data <= 8'hF8;
            16'd3298: data <= 8'h00;
            16'd3299: data <= 8'hF8;
            16'd3300: data <= 8'h00;
            16'd3301: data <= 8'hF8;
            16'd3302: data <= 8'h00;
            16'd3303: data <= 8'hF8;
            16'd3304: data <= 8'h00;
            16'd3305: data <= 8'hF8;
            16'd3306: data <= 8'h00;
            16'd3307: data <= 8'hF8;
            16'd3308: data <= 8'h00;
            16'd3309: data <= 8'hF8;
            16'd3310: data <= 8'h00;
            16'd3311: data <= 8'hF8;
            16'd3312: data <= 8'h00;
            16'd3313: data <= 8'hF8;
            16'd3314: data <= 8'h00;
            16'd3315: data <= 8'hF8;
            16'd3316: data <= 8'h00;
            16'd3317: data <= 8'hF8;
            16'd3318: data <= 8'h00;
            16'd3319: data <= 8'hF8;
            16'd3320: data <= 8'hFF;
            16'd3321: data <= 8'hFF;
            16'd3322: data <= 8'h00;
            16'd3323: data <= 8'hF8;
            16'd3324: data <= 8'h00;
            16'd3325: data <= 8'hF8;
            16'd3326: data <= 8'h00;
            16'd3327: data <= 8'hF8;
            16'd3328: data <= 8'h00;
            16'd3329: data <= 8'hF8;
            16'd3330: data <= 8'h00;
            16'd3331: data <= 8'hF8;
            16'd3332: data <= 8'h00;
            16'd3333: data <= 8'hF8;
            16'd3334: data <= 8'h00;
            16'd3335: data <= 8'hF8;
            16'd3336: data <= 8'h00;
            16'd3337: data <= 8'hF8;
            16'd3338: data <= 8'h00;
            16'd3339: data <= 8'hF8;
            16'd3340: data <= 8'h00;
            16'd3341: data <= 8'hF8;
            16'd3342: data <= 8'h00;
            16'd3343: data <= 8'hF8;
            16'd3344: data <= 8'h00;
            16'd3345: data <= 8'hF8;
            16'd3346: data <= 8'h00;
            16'd3347: data <= 8'hF8;
            16'd3348: data <= 8'h00;
            16'd3349: data <= 8'hF8;
            16'd3350: data <= 8'h00;
            16'd3351: data <= 8'hF8;
            16'd3352: data <= 8'h00;
            16'd3353: data <= 8'hF8;
            16'd3354: data <= 8'h00;
            16'd3355: data <= 8'hF8;
            16'd3356: data <= 8'h00;
            16'd3357: data <= 8'hF8;
            16'd3358: data <= 8'h00;
            16'd3359: data <= 8'hF8;
            16'd3360: data <= 8'hFF;
            16'd3361: data <= 8'hFF;
            16'd3362: data <= 8'h00;
            16'd3363: data <= 8'hF8;
            16'd3364: data <= 8'h00;
            16'd3365: data <= 8'hF8;
            16'd3366: data <= 8'h00;
            16'd3367: data <= 8'hF8;
            16'd3368: data <= 8'h00;
            16'd3369: data <= 8'hF8;
            16'd3370: data <= 8'h00;
            16'd3371: data <= 8'hF8;
            16'd3372: data <= 8'h00;
            16'd3373: data <= 8'hF8;
            16'd3374: data <= 8'h00;
            16'd3375: data <= 8'hF8;
            16'd3376: data <= 8'h00;
            16'd3377: data <= 8'hF8;
            16'd3378: data <= 8'h00;
            16'd3379: data <= 8'hF8;
            16'd3380: data <= 8'h00;
            16'd3381: data <= 8'hF8;
            16'd3382: data <= 8'h00;
            16'd3383: data <= 8'hF8;
            16'd3384: data <= 8'h00;
            16'd3385: data <= 8'hF8;
            16'd3386: data <= 8'h00;
            16'd3387: data <= 8'hF8;
            16'd3388: data <= 8'h00;
            16'd3389: data <= 8'hF8;
            16'd3390: data <= 8'h00;
            16'd3391: data <= 8'hF8;
            16'd3392: data <= 8'h00;
            16'd3393: data <= 8'hF8;
            16'd3394: data <= 8'h00;
            16'd3395: data <= 8'hF8;
            16'd3396: data <= 8'h00;
            16'd3397: data <= 8'hF8;
            16'd3398: data <= 8'h00;
            16'd3399: data <= 8'hF8;
            16'd3400: data <= 8'hFF;
            16'd3401: data <= 8'hFF;
            16'd3402: data <= 8'h00;
            16'd3403: data <= 8'hF8;
            16'd3404: data <= 8'h00;
            16'd3405: data <= 8'hF8;
            16'd3406: data <= 8'h00;
            16'd3407: data <= 8'hF8;
            16'd3408: data <= 8'h00;
            16'd3409: data <= 8'hF8;
            16'd3410: data <= 8'h00;
            16'd3411: data <= 8'hF8;
            16'd3412: data <= 8'h00;
            16'd3413: data <= 8'hF8;
            16'd3414: data <= 8'h00;
            16'd3415: data <= 8'hF8;
            16'd3416: data <= 8'h00;
            16'd3417: data <= 8'hF8;
            16'd3418: data <= 8'h00;
            16'd3419: data <= 8'hF8;
            16'd3420: data <= 8'h00;
            16'd3421: data <= 8'hF8;
            16'd3422: data <= 8'h00;
            16'd3423: data <= 8'hF8;
            16'd3424: data <= 8'h00;
            16'd3425: data <= 8'hF8;
            16'd3426: data <= 8'h00;
            16'd3427: data <= 8'hF8;
            16'd3428: data <= 8'h00;
            16'd3429: data <= 8'hF8;
            16'd3430: data <= 8'h00;
            16'd3431: data <= 8'hF8;
            16'd3432: data <= 8'h00;
            16'd3433: data <= 8'hF8;
            16'd3434: data <= 8'h00;
            16'd3435: data <= 8'hF8;
            16'd3436: data <= 8'h00;
            16'd3437: data <= 8'hF8;
            16'd3438: data <= 8'h00;
            16'd3439: data <= 8'hF8;
            16'd3440: data <= 8'hFF;
            16'd3441: data <= 8'hFF;
            16'd3442: data <= 8'h00;
            16'd3443: data <= 8'hF8;
            16'd3444: data <= 8'h00;
            16'd3445: data <= 8'hF8;
            16'd3446: data <= 8'h00;
            16'd3447: data <= 8'hF8;
            16'd3448: data <= 8'h00;
            16'd3449: data <= 8'hF8;
            16'd3450: data <= 8'h00;
            16'd3451: data <= 8'hF8;
            16'd3452: data <= 8'h00;
            16'd3453: data <= 8'hF8;
            16'd3454: data <= 8'h00;
            16'd3455: data <= 8'hF8;
            16'd3456: data <= 8'h00;
            16'd3457: data <= 8'hF8;
            16'd3458: data <= 8'h00;
            16'd3459: data <= 8'hF8;
            16'd3460: data <= 8'h00;
            16'd3461: data <= 8'hF8;
            16'd3462: data <= 8'h00;
            16'd3463: data <= 8'hF8;
            16'd3464: data <= 8'h00;
            16'd3465: data <= 8'hF8;
            16'd3466: data <= 8'h00;
            16'd3467: data <= 8'hF8;
            16'd3468: data <= 8'h00;
            16'd3469: data <= 8'hF8;
            16'd3470: data <= 8'h00;
            16'd3471: data <= 8'hF8;
            16'd3472: data <= 8'h00;
            16'd3473: data <= 8'hF8;
            16'd3474: data <= 8'h00;
            16'd3475: data <= 8'hF8;
            16'd3476: data <= 8'h00;
            16'd3477: data <= 8'hF8;
            16'd3478: data <= 8'h00;
            16'd3479: data <= 8'hF8;
            16'd3480: data <= 8'hFF;
            16'd3481: data <= 8'hFF;
            16'd3482: data <= 8'h00;
            16'd3483: data <= 8'hF8;
            16'd3484: data <= 8'h00;
            16'd3485: data <= 8'hF8;
            16'd3486: data <= 8'h00;
            16'd3487: data <= 8'hF8;
            16'd3488: data <= 8'h00;
            16'd3489: data <= 8'hF8;
            16'd3490: data <= 8'h00;
            16'd3491: data <= 8'hF8;
            16'd3492: data <= 8'h00;
            16'd3493: data <= 8'hF8;
            16'd3494: data <= 8'h00;
            16'd3495: data <= 8'hF8;
            16'd3496: data <= 8'h00;
            16'd3497: data <= 8'hF8;
            16'd3498: data <= 8'h00;
            16'd3499: data <= 8'hF8;
            16'd3500: data <= 8'h00;
            16'd3501: data <= 8'hF8;
            16'd3502: data <= 8'h00;
            16'd3503: data <= 8'hF8;
            16'd3504: data <= 8'h00;
            16'd3505: data <= 8'hF8;
            16'd3506: data <= 8'h00;
            16'd3507: data <= 8'hF8;
            16'd3508: data <= 8'h00;
            16'd3509: data <= 8'hF8;
            16'd3510: data <= 8'h00;
            16'd3511: data <= 8'hF8;
            16'd3512: data <= 8'h00;
            16'd3513: data <= 8'hF8;
            16'd3514: data <= 8'h00;
            16'd3515: data <= 8'hF8;
            16'd3516: data <= 8'h00;
            16'd3517: data <= 8'hF8;
            16'd3518: data <= 8'h00;
            16'd3519: data <= 8'hF8;
            16'd3520: data <= 8'hFF;
            16'd3521: data <= 8'hFF;
            16'd3522: data <= 8'h00;
            16'd3523: data <= 8'hF8;
            16'd3524: data <= 8'h00;
            16'd3525: data <= 8'hF8;
            16'd3526: data <= 8'h00;
            16'd3527: data <= 8'hF8;
            16'd3528: data <= 8'h00;
            16'd3529: data <= 8'hF8;
            16'd3530: data <= 8'h00;
            16'd3531: data <= 8'hF8;
            16'd3532: data <= 8'h00;
            16'd3533: data <= 8'hF8;
            16'd3534: data <= 8'h00;
            16'd3535: data <= 8'hF8;
            16'd3536: data <= 8'h00;
            16'd3537: data <= 8'hF8;
            16'd3538: data <= 8'h00;
            16'd3539: data <= 8'hF8;
            16'd3540: data <= 8'h00;
            16'd3541: data <= 8'hF8;
            16'd3542: data <= 8'h00;
            16'd3543: data <= 8'hF8;
            16'd3544: data <= 8'h00;
            16'd3545: data <= 8'hF8;
            16'd3546: data <= 8'h00;
            16'd3547: data <= 8'hF8;
            16'd3548: data <= 8'h00;
            16'd3549: data <= 8'hF8;
            16'd3550: data <= 8'h00;
            16'd3551: data <= 8'hF8;
            16'd3552: data <= 8'h00;
            16'd3553: data <= 8'hF8;
            16'd3554: data <= 8'h00;
            16'd3555: data <= 8'hF8;
            16'd3556: data <= 8'h00;
            16'd3557: data <= 8'hF8;
            16'd3558: data <= 8'h00;
            16'd3559: data <= 8'hF8;
            16'd3560: data <= 8'hFF;
            16'd3561: data <= 8'hFF;
            16'd3562: data <= 8'h00;
            16'd3563: data <= 8'hF8;
            16'd3564: data <= 8'h00;
            16'd3565: data <= 8'hF8;
            16'd3566: data <= 8'h00;
            16'd3567: data <= 8'hF8;
            16'd3568: data <= 8'h00;
            16'd3569: data <= 8'hF8;
            16'd3570: data <= 8'h00;
            16'd3571: data <= 8'hF8;
            16'd3572: data <= 8'h00;
            16'd3573: data <= 8'hF8;
            16'd3574: data <= 8'h00;
            16'd3575: data <= 8'hF8;
            16'd3576: data <= 8'h00;
            16'd3577: data <= 8'hF8;
            16'd3578: data <= 8'h00;
            16'd3579: data <= 8'hF8;
            16'd3580: data <= 8'h00;
            16'd3581: data <= 8'hF8;
            16'd3582: data <= 8'h00;
            16'd3583: data <= 8'hF8;
            16'd3584: data <= 8'h00;
            16'd3585: data <= 8'hF8;
            16'd3586: data <= 8'h00;
            16'd3587: data <= 8'hF8;
            16'd3588: data <= 8'h00;
            16'd3589: data <= 8'hF8;
            16'd3590: data <= 8'h00;
            16'd3591: data <= 8'hF8;
            16'd3592: data <= 8'h00;
            16'd3593: data <= 8'hF8;
            16'd3594: data <= 8'h00;
            16'd3595: data <= 8'hF8;
            16'd3596: data <= 8'h00;
            16'd3597: data <= 8'hF8;
            16'd3598: data <= 8'h00;
            16'd3599: data <= 8'hF8;
            16'd3600: data <= 8'hFF;
            16'd3601: data <= 8'hFF;
            16'd3602: data <= 8'h00;
            16'd3603: data <= 8'hF8;
            16'd3604: data <= 8'h00;
            16'd3605: data <= 8'hF8;
            16'd3606: data <= 8'h00;
            16'd3607: data <= 8'hF8;
            16'd3608: data <= 8'h00;
            16'd3609: data <= 8'hF8;
            16'd3610: data <= 8'h00;
            16'd3611: data <= 8'hF8;
            16'd3612: data <= 8'h00;
            16'd3613: data <= 8'hF8;
            16'd3614: data <= 8'h00;
            16'd3615: data <= 8'hF8;
            16'd3616: data <= 8'h00;
            16'd3617: data <= 8'hF8;
            16'd3618: data <= 8'h00;
            16'd3619: data <= 8'hF8;
            16'd3620: data <= 8'h00;
            16'd3621: data <= 8'hF8;
            16'd3622: data <= 8'h00;
            16'd3623: data <= 8'hF8;
            16'd3624: data <= 8'h00;
            16'd3625: data <= 8'hF8;
            16'd3626: data <= 8'h00;
            16'd3627: data <= 8'hF8;
            16'd3628: data <= 8'h00;
            16'd3629: data <= 8'hF8;
            16'd3630: data <= 8'h00;
            16'd3631: data <= 8'hF8;
            16'd3632: data <= 8'h00;
            16'd3633: data <= 8'hF8;
            16'd3634: data <= 8'h00;
            16'd3635: data <= 8'hF8;
            16'd3636: data <= 8'h00;
            16'd3637: data <= 8'hF8;
            16'd3638: data <= 8'h00;
            16'd3639: data <= 8'hF8;
            16'd3640: data <= 8'hFF;
            16'd3641: data <= 8'hFF;
            16'd3642: data <= 8'h00;
            16'd3643: data <= 8'hF8;
            16'd3644: data <= 8'h00;
            16'd3645: data <= 8'hF8;
            16'd3646: data <= 8'h00;
            16'd3647: data <= 8'hF8;
            16'd3648: data <= 8'h00;
            16'd3649: data <= 8'hF8;
            16'd3650: data <= 8'h00;
            16'd3651: data <= 8'hF8;
            16'd3652: data <= 8'h00;
            16'd3653: data <= 8'hF8;
            16'd3654: data <= 8'h00;
            16'd3655: data <= 8'hF8;
            16'd3656: data <= 8'h00;
            16'd3657: data <= 8'hF8;
            16'd3658: data <= 8'h00;
            16'd3659: data <= 8'hF8;
            16'd3660: data <= 8'h00;
            16'd3661: data <= 8'hF8;
            16'd3662: data <= 8'h00;
            16'd3663: data <= 8'hF8;
            16'd3664: data <= 8'h00;
            16'd3665: data <= 8'hF8;
            16'd3666: data <= 8'h00;
            16'd3667: data <= 8'hF8;
            16'd3668: data <= 8'h00;
            16'd3669: data <= 8'hF8;
            16'd3670: data <= 8'h00;
            16'd3671: data <= 8'hF8;
            16'd3672: data <= 8'h00;
            16'd3673: data <= 8'hF8;
            16'd3674: data <= 8'h00;
            16'd3675: data <= 8'hF8;
            16'd3676: data <= 8'h00;
            16'd3677: data <= 8'hF8;
            16'd3678: data <= 8'h00;
            16'd3679: data <= 8'hF8;
            16'd3680: data <= 8'hFF;
            16'd3681: data <= 8'hFF;
            16'd3682: data <= 8'h00;
            16'd3683: data <= 8'hF8;
            16'd3684: data <= 8'h00;
            16'd3685: data <= 8'hF8;
            16'd3686: data <= 8'h00;
            16'd3687: data <= 8'hF8;
            16'd3688: data <= 8'h00;
            16'd3689: data <= 8'hF8;
            16'd3690: data <= 8'h00;
            16'd3691: data <= 8'hF8;
            16'd3692: data <= 8'h00;
            16'd3693: data <= 8'hF8;
            16'd3694: data <= 8'h00;
            16'd3695: data <= 8'hF8;
            16'd3696: data <= 8'h00;
            16'd3697: data <= 8'hF8;
            16'd3698: data <= 8'h00;
            16'd3699: data <= 8'hF8;
            16'd3700: data <= 8'h00;
            16'd3701: data <= 8'hF8;
            16'd3702: data <= 8'h00;
            16'd3703: data <= 8'hF8;
            16'd3704: data <= 8'h00;
            16'd3705: data <= 8'hF8;
            16'd3706: data <= 8'h00;
            16'd3707: data <= 8'hF8;
            16'd3708: data <= 8'h00;
            16'd3709: data <= 8'hF8;
            16'd3710: data <= 8'h00;
            16'd3711: data <= 8'hF8;
            16'd3712: data <= 8'h00;
            16'd3713: data <= 8'hF8;
            16'd3714: data <= 8'h00;
            16'd3715: data <= 8'hF8;
            16'd3716: data <= 8'h00;
            16'd3717: data <= 8'hF8;
            16'd3718: data <= 8'h00;
            16'd3719: data <= 8'hF8;
            16'd3720: data <= 8'hFF;
            16'd3721: data <= 8'hFF;
            16'd3722: data <= 8'h00;
            16'd3723: data <= 8'hF8;
            16'd3724: data <= 8'h00;
            16'd3725: data <= 8'hF8;
            16'd3726: data <= 8'h00;
            16'd3727: data <= 8'hF8;
            16'd3728: data <= 8'h00;
            16'd3729: data <= 8'hF8;
            16'd3730: data <= 8'h00;
            16'd3731: data <= 8'hF8;
            16'd3732: data <= 8'h00;
            16'd3733: data <= 8'hF8;
            16'd3734: data <= 8'h00;
            16'd3735: data <= 8'hF8;
            16'd3736: data <= 8'h00;
            16'd3737: data <= 8'hF8;
            16'd3738: data <= 8'h00;
            16'd3739: data <= 8'hF8;
            16'd3740: data <= 8'h00;
            16'd3741: data <= 8'hF8;
            16'd3742: data <= 8'h00;
            16'd3743: data <= 8'hF8;
            16'd3744: data <= 8'h00;
            16'd3745: data <= 8'hF8;
            16'd3746: data <= 8'h00;
            16'd3747: data <= 8'hF8;
            16'd3748: data <= 8'h00;
            16'd3749: data <= 8'hF8;
            16'd3750: data <= 8'h00;
            16'd3751: data <= 8'hF8;
            16'd3752: data <= 8'h00;
            16'd3753: data <= 8'hF8;
            16'd3754: data <= 8'h00;
            16'd3755: data <= 8'hF8;
            16'd3756: data <= 8'h00;
            16'd3757: data <= 8'hF8;
            16'd3758: data <= 8'h00;
            16'd3759: data <= 8'hF8;
            16'd3760: data <= 8'hFF;
            16'd3761: data <= 8'hFF;
            16'd3762: data <= 8'h00;
            16'd3763: data <= 8'hF8;
            16'd3764: data <= 8'h00;
            16'd3765: data <= 8'hF8;
            16'd3766: data <= 8'h00;
            16'd3767: data <= 8'hF8;
            16'd3768: data <= 8'h00;
            16'd3769: data <= 8'hF8;
            16'd3770: data <= 8'h00;
            16'd3771: data <= 8'hF8;
            16'd3772: data <= 8'h00;
            16'd3773: data <= 8'hF8;
            16'd3774: data <= 8'h00;
            16'd3775: data <= 8'hF8;
            16'd3776: data <= 8'h00;
            16'd3777: data <= 8'hF8;
            16'd3778: data <= 8'h00;
            16'd3779: data <= 8'hF8;
            16'd3780: data <= 8'h00;
            16'd3781: data <= 8'hF8;
            16'd3782: data <= 8'h00;
            16'd3783: data <= 8'hF8;
            16'd3784: data <= 8'h00;
            16'd3785: data <= 8'hF8;
            16'd3786: data <= 8'h00;
            16'd3787: data <= 8'hF8;
            16'd3788: data <= 8'h00;
            16'd3789: data <= 8'hF8;
            16'd3790: data <= 8'h00;
            16'd3791: data <= 8'hF8;
            16'd3792: data <= 8'h00;
            16'd3793: data <= 8'hF8;
            16'd3794: data <= 8'h00;
            16'd3795: data <= 8'hF8;
            16'd3796: data <= 8'h00;
            16'd3797: data <= 8'hF8;
            16'd3798: data <= 8'h00;
            16'd3799: data <= 8'hF8;
            16'd3800: data <= 8'hFF;
            16'd3801: data <= 8'hFF;
            16'd3802: data <= 8'h00;
            16'd3803: data <= 8'hF8;
            16'd3804: data <= 8'h00;
            16'd3805: data <= 8'hF8;
            16'd3806: data <= 8'h00;
            16'd3807: data <= 8'hF8;
            16'd3808: data <= 8'h00;
            16'd3809: data <= 8'hF8;
            16'd3810: data <= 8'h00;
            16'd3811: data <= 8'hF8;
            16'd3812: data <= 8'h00;
            16'd3813: data <= 8'hF8;
            16'd3814: data <= 8'h00;
            16'd3815: data <= 8'hF8;
            16'd3816: data <= 8'h00;
            16'd3817: data <= 8'hF8;
            16'd3818: data <= 8'h00;
            16'd3819: data <= 8'hF8;
            16'd3820: data <= 8'h00;
            16'd3821: data <= 8'hF8;
            16'd3822: data <= 8'h00;
            16'd3823: data <= 8'hF8;
            16'd3824: data <= 8'h00;
            16'd3825: data <= 8'hF8;
            16'd3826: data <= 8'h00;
            16'd3827: data <= 8'hF8;
            16'd3828: data <= 8'h00;
            16'd3829: data <= 8'hF8;
            16'd3830: data <= 8'h00;
            16'd3831: data <= 8'hF8;
            16'd3832: data <= 8'h00;
            16'd3833: data <= 8'hF8;
            16'd3834: data <= 8'h00;
            16'd3835: data <= 8'hF8;
            16'd3836: data <= 8'h00;
            16'd3837: data <= 8'hF8;
            16'd3838: data <= 8'h00;
            16'd3839: data <= 8'hF8;
            16'd3840: data <= 8'hFF;
            16'd3841: data <= 8'hFF;
            16'd3842: data <= 8'h00;
            16'd3843: data <= 8'hF8;
            16'd3844: data <= 8'h00;
            16'd3845: data <= 8'hF8;
            16'd3846: data <= 8'h00;
            16'd3847: data <= 8'hF8;
            16'd3848: data <= 8'h00;
            16'd3849: data <= 8'hF8;
            16'd3850: data <= 8'h00;
            16'd3851: data <= 8'hF8;
            16'd3852: data <= 8'h00;
            16'd3853: data <= 8'hF8;
            16'd3854: data <= 8'h00;
            16'd3855: data <= 8'hF8;
            16'd3856: data <= 8'h00;
            16'd3857: data <= 8'hF8;
            16'd3858: data <= 8'h00;
            16'd3859: data <= 8'hF8;
            16'd3860: data <= 8'h00;
            16'd3861: data <= 8'hF8;
            16'd3862: data <= 8'h00;
            16'd3863: data <= 8'hF8;
            16'd3864: data <= 8'h00;
            16'd3865: data <= 8'hF8;
            16'd3866: data <= 8'h00;
            16'd3867: data <= 8'hF8;
            16'd3868: data <= 8'h00;
            16'd3869: data <= 8'hF8;
            16'd3870: data <= 8'h00;
            16'd3871: data <= 8'hF8;
            16'd3872: data <= 8'h00;
            16'd3873: data <= 8'hF8;
            16'd3874: data <= 8'h00;
            16'd3875: data <= 8'hF8;
            16'd3876: data <= 8'h00;
            16'd3877: data <= 8'hF8;
            16'd3878: data <= 8'h00;
            16'd3879: data <= 8'hF8;
            16'd3880: data <= 8'hFF;
            16'd3881: data <= 8'hFF;
            16'd3882: data <= 8'h00;
            16'd3883: data <= 8'hF8;
            16'd3884: data <= 8'h00;
            16'd3885: data <= 8'hF8;
            16'd3886: data <= 8'h00;
            16'd3887: data <= 8'hF8;
            16'd3888: data <= 8'h00;
            16'd3889: data <= 8'hF8;
            16'd3890: data <= 8'h00;
            16'd3891: data <= 8'hF8;
            16'd3892: data <= 8'h00;
            16'd3893: data <= 8'hF8;
            16'd3894: data <= 8'h00;
            16'd3895: data <= 8'hF8;
            16'd3896: data <= 8'h00;
            16'd3897: data <= 8'hF8;
            16'd3898: data <= 8'h00;
            16'd3899: data <= 8'hF8;
            16'd3900: data <= 8'h00;
            16'd3901: data <= 8'hF8;
            16'd3902: data <= 8'h00;
            16'd3903: data <= 8'hF8;
            16'd3904: data <= 8'h00;
            16'd3905: data <= 8'hF8;
            16'd3906: data <= 8'h00;
            16'd3907: data <= 8'hF8;
            16'd3908: data <= 8'h00;
            16'd3909: data <= 8'hF8;
            16'd3910: data <= 8'h00;
            16'd3911: data <= 8'hF8;
            16'd3912: data <= 8'h00;
            16'd3913: data <= 8'hF8;
            16'd3914: data <= 8'h00;
            16'd3915: data <= 8'hF8;
            16'd3916: data <= 8'h00;
            16'd3917: data <= 8'hF8;
            16'd3918: data <= 8'h00;
            16'd3919: data <= 8'hF8;
            16'd3920: data <= 8'hFF;
            16'd3921: data <= 8'hFF;
            16'd3922: data <= 8'h00;
            16'd3923: data <= 8'hF8;
            16'd3924: data <= 8'h00;
            16'd3925: data <= 8'hF8;
            16'd3926: data <= 8'h00;
            16'd3927: data <= 8'hF8;
            16'd3928: data <= 8'h00;
            16'd3929: data <= 8'hF8;
            16'd3930: data <= 8'h00;
            16'd3931: data <= 8'hF8;
            16'd3932: data <= 8'h00;
            16'd3933: data <= 8'hF8;
            16'd3934: data <= 8'h00;
            16'd3935: data <= 8'hF8;
            16'd3936: data <= 8'h00;
            16'd3937: data <= 8'hF8;
            16'd3938: data <= 8'h00;
            16'd3939: data <= 8'hF8;
            16'd3940: data <= 8'h00;
            16'd3941: data <= 8'hF8;
            16'd3942: data <= 8'h00;
            16'd3943: data <= 8'hF8;
            16'd3944: data <= 8'h00;
            16'd3945: data <= 8'hF8;
            16'd3946: data <= 8'h00;
            16'd3947: data <= 8'hF8;
            16'd3948: data <= 8'h00;
            16'd3949: data <= 8'hF8;
            16'd3950: data <= 8'h00;
            16'd3951: data <= 8'hF8;
            16'd3952: data <= 8'h00;
            16'd3953: data <= 8'hF8;
            16'd3954: data <= 8'h00;
            16'd3955: data <= 8'hF8;
            16'd3956: data <= 8'h00;
            16'd3957: data <= 8'hF8;
            16'd3958: data <= 8'h00;
            16'd3959: data <= 8'hF8;
            16'd3960: data <= 8'hFF;
            16'd3961: data <= 8'hFF;
            16'd3962: data <= 8'h00;
            16'd3963: data <= 8'hF8;
            16'd3964: data <= 8'h00;
            16'd3965: data <= 8'hF8;
            16'd3966: data <= 8'h00;
            16'd3967: data <= 8'hF8;
            16'd3968: data <= 8'h00;
            16'd3969: data <= 8'hF8;
            16'd3970: data <= 8'h00;
            16'd3971: data <= 8'hF8;
            16'd3972: data <= 8'h00;
            16'd3973: data <= 8'hF8;
            16'd3974: data <= 8'h00;
            16'd3975: data <= 8'hF8;
            16'd3976: data <= 8'h00;
            16'd3977: data <= 8'hF8;
            16'd3978: data <= 8'h00;
            16'd3979: data <= 8'hF8;
            16'd3980: data <= 8'h00;
            16'd3981: data <= 8'hF8;
            16'd3982: data <= 8'h00;
            16'd3983: data <= 8'hF8;
            16'd3984: data <= 8'h00;
            16'd3985: data <= 8'hF8;
            16'd3986: data <= 8'h00;
            16'd3987: data <= 8'hF8;
            16'd3988: data <= 8'h00;
            16'd3989: data <= 8'hF8;
            16'd3990: data <= 8'h00;
            16'd3991: data <= 8'hF8;
            16'd3992: data <= 8'h00;
            16'd3993: data <= 8'hF8;
            16'd3994: data <= 8'h00;
            16'd3995: data <= 8'hF8;
            16'd3996: data <= 8'h00;
            16'd3997: data <= 8'hF8;
            16'd3998: data <= 8'h00;
            16'd3999: data <= 8'hF8;
            16'd4000: data <= 8'hFF;
            16'd4001: data <= 8'hFF;
            16'd4002: data <= 8'h00;
            16'd4003: data <= 8'hF8;
            16'd4004: data <= 8'h00;
            16'd4005: data <= 8'hF8;
            16'd4006: data <= 8'h00;
            16'd4007: data <= 8'hF8;
            16'd4008: data <= 8'h00;
            16'd4009: data <= 8'hF8;
            16'd4010: data <= 8'h00;
            16'd4011: data <= 8'hF8;
            16'd4012: data <= 8'h00;
            16'd4013: data <= 8'hF8;
            16'd4014: data <= 8'h00;
            16'd4015: data <= 8'hF8;
            16'd4016: data <= 8'h00;
            16'd4017: data <= 8'hF8;
            16'd4018: data <= 8'h00;
            16'd4019: data <= 8'hF8;
            16'd4020: data <= 8'h00;
            16'd4021: data <= 8'hF8;
            16'd4022: data <= 8'h00;
            16'd4023: data <= 8'hF8;
            16'd4024: data <= 8'h00;
            16'd4025: data <= 8'hF8;
            16'd4026: data <= 8'h00;
            16'd4027: data <= 8'hF8;
            16'd4028: data <= 8'h00;
            16'd4029: data <= 8'hF8;
            16'd4030: data <= 8'h00;
            16'd4031: data <= 8'hF8;
            16'd4032: data <= 8'h00;
            16'd4033: data <= 8'hF8;
            16'd4034: data <= 8'h00;
            16'd4035: data <= 8'hF8;
            16'd4036: data <= 8'h00;
            16'd4037: data <= 8'hF8;
            16'd4038: data <= 8'h00;
            16'd4039: data <= 8'hF8;
            16'd4040: data <= 8'hFF;
            16'd4041: data <= 8'hFF;
            16'd4042: data <= 8'h00;
            16'd4043: data <= 8'hF8;
            16'd4044: data <= 8'h00;
            16'd4045: data <= 8'hF8;
            16'd4046: data <= 8'h00;
            16'd4047: data <= 8'hF8;
            16'd4048: data <= 8'h00;
            16'd4049: data <= 8'hF8;
            16'd4050: data <= 8'h00;
            16'd4051: data <= 8'hF8;
            16'd4052: data <= 8'h00;
            16'd4053: data <= 8'hF8;
            16'd4054: data <= 8'h00;
            16'd4055: data <= 8'hF8;
            16'd4056: data <= 8'h00;
            16'd4057: data <= 8'hF8;
            16'd4058: data <= 8'h00;
            16'd4059: data <= 8'hF8;
            16'd4060: data <= 8'h00;
            16'd4061: data <= 8'hF8;
            16'd4062: data <= 8'h00;
            16'd4063: data <= 8'hF8;
            16'd4064: data <= 8'h00;
            16'd4065: data <= 8'hF8;
            16'd4066: data <= 8'h00;
            16'd4067: data <= 8'hF8;
            16'd4068: data <= 8'h00;
            16'd4069: data <= 8'hF8;
            16'd4070: data <= 8'h00;
            16'd4071: data <= 8'hF8;
            16'd4072: data <= 8'h00;
            16'd4073: data <= 8'hF8;
            16'd4074: data <= 8'h00;
            16'd4075: data <= 8'hF8;
            16'd4076: data <= 8'h00;
            16'd4077: data <= 8'hF8;
            16'd4078: data <= 8'h00;
            16'd4079: data <= 8'hF8;
            16'd4080: data <= 8'hFF;
            16'd4081: data <= 8'hFF;
            16'd4082: data <= 8'h00;
            16'd4083: data <= 8'hF8;
            16'd4084: data <= 8'h00;
            16'd4085: data <= 8'hF8;
            16'd4086: data <= 8'h00;
            16'd4087: data <= 8'hF8;
            16'd4088: data <= 8'h00;
            16'd4089: data <= 8'hF8;
            16'd4090: data <= 8'h00;
            16'd4091: data <= 8'hF8;
            16'd4092: data <= 8'h00;
            16'd4093: data <= 8'hF8;
            16'd4094: data <= 8'h00;
            16'd4095: data <= 8'hF8;
            16'd4096: data <= 8'h00;
            16'd4097: data <= 8'hF8;
            16'd4098: data <= 8'h00;
            16'd4099: data <= 8'hF8;
            16'd4100: data <= 8'h00;
            16'd4101: data <= 8'hF8;
            16'd4102: data <= 8'h00;
            16'd4103: data <= 8'hF8;
            16'd4104: data <= 8'h00;
            16'd4105: data <= 8'hF8;
            16'd4106: data <= 8'h00;
            16'd4107: data <= 8'hF8;
            16'd4108: data <= 8'h00;
            16'd4109: data <= 8'hF8;
            16'd4110: data <= 8'h00;
            16'd4111: data <= 8'hF8;
            16'd4112: data <= 8'h00;
            16'd4113: data <= 8'hF8;
            16'd4114: data <= 8'h00;
            16'd4115: data <= 8'hF8;
            16'd4116: data <= 8'h00;
            16'd4117: data <= 8'hF8;
            16'd4118: data <= 8'h00;
            16'd4119: data <= 8'hF8;
            16'd4120: data <= 8'hFF;
            16'd4121: data <= 8'hFF;
            16'd4122: data <= 8'h00;
            16'd4123: data <= 8'hF8;
            16'd4124: data <= 8'h00;
            16'd4125: data <= 8'hF8;
            16'd4126: data <= 8'h00;
            16'd4127: data <= 8'hF8;
            16'd4128: data <= 8'h00;
            16'd4129: data <= 8'hF8;
            16'd4130: data <= 8'h00;
            16'd4131: data <= 8'hF8;
            16'd4132: data <= 8'h00;
            16'd4133: data <= 8'hF8;
            16'd4134: data <= 8'h00;
            16'd4135: data <= 8'hF8;
            16'd4136: data <= 8'h00;
            16'd4137: data <= 8'hF8;
            16'd4138: data <= 8'h00;
            16'd4139: data <= 8'hF8;
            16'd4140: data <= 8'h00;
            16'd4141: data <= 8'hF8;
            16'd4142: data <= 8'h00;
            16'd4143: data <= 8'hF8;
            16'd4144: data <= 8'h00;
            16'd4145: data <= 8'hF8;
            16'd4146: data <= 8'h00;
            16'd4147: data <= 8'hF8;
            16'd4148: data <= 8'h00;
            16'd4149: data <= 8'hF8;
            16'd4150: data <= 8'h00;
            16'd4151: data <= 8'hF8;
            16'd4152: data <= 8'h00;
            16'd4153: data <= 8'hF8;
            16'd4154: data <= 8'h00;
            16'd4155: data <= 8'hF8;
            16'd4156: data <= 8'h00;
            16'd4157: data <= 8'hF8;
            16'd4158: data <= 8'h00;
            16'd4159: data <= 8'hF8;
            16'd4160: data <= 8'hFF;
            16'd4161: data <= 8'hFF;
            16'd4162: data <= 8'h00;
            16'd4163: data <= 8'hF8;
            16'd4164: data <= 8'h00;
            16'd4165: data <= 8'hF8;
            16'd4166: data <= 8'h00;
            16'd4167: data <= 8'hF8;
            16'd4168: data <= 8'h00;
            16'd4169: data <= 8'hF8;
            16'd4170: data <= 8'h00;
            16'd4171: data <= 8'hF8;
            16'd4172: data <= 8'h00;
            16'd4173: data <= 8'hF8;
            16'd4174: data <= 8'h00;
            16'd4175: data <= 8'hF8;
            16'd4176: data <= 8'h00;
            16'd4177: data <= 8'hF8;
            16'd4178: data <= 8'h00;
            16'd4179: data <= 8'hF8;
            16'd4180: data <= 8'h00;
            16'd4181: data <= 8'hF8;
            16'd4182: data <= 8'h00;
            16'd4183: data <= 8'hF8;
            16'd4184: data <= 8'h00;
            16'd4185: data <= 8'hF8;
            16'd4186: data <= 8'h00;
            16'd4187: data <= 8'hF8;
            16'd4188: data <= 8'h00;
            16'd4189: data <= 8'hF8;
            16'd4190: data <= 8'h00;
            16'd4191: data <= 8'hF8;
            16'd4192: data <= 8'h00;
            16'd4193: data <= 8'hF8;
            16'd4194: data <= 8'h00;
            16'd4195: data <= 8'hF8;
            16'd4196: data <= 8'h00;
            16'd4197: data <= 8'hF8;
            16'd4198: data <= 8'h00;
            16'd4199: data <= 8'hF8;
            16'd4200: data <= 8'hFF;
            16'd4201: data <= 8'hFF;
            16'd4202: data <= 8'h00;
            16'd4203: data <= 8'hF8;
            16'd4204: data <= 8'h00;
            16'd4205: data <= 8'hF8;
            16'd4206: data <= 8'h00;
            16'd4207: data <= 8'hF8;
            16'd4208: data <= 8'h00;
            16'd4209: data <= 8'hF8;
            16'd4210: data <= 8'h00;
            16'd4211: data <= 8'hF8;
            16'd4212: data <= 8'h00;
            16'd4213: data <= 8'hF8;
            16'd4214: data <= 8'h00;
            16'd4215: data <= 8'hF8;
            16'd4216: data <= 8'h00;
            16'd4217: data <= 8'hF8;
            16'd4218: data <= 8'h00;
            16'd4219: data <= 8'hF8;
            16'd4220: data <= 8'h00;
            16'd4221: data <= 8'hF8;
            16'd4222: data <= 8'h00;
            16'd4223: data <= 8'hF8;
            16'd4224: data <= 8'h00;
            16'd4225: data <= 8'hF8;
            16'd4226: data <= 8'h00;
            16'd4227: data <= 8'hF8;
            16'd4228: data <= 8'h00;
            16'd4229: data <= 8'hF8;
            16'd4230: data <= 8'h00;
            16'd4231: data <= 8'hF8;
            16'd4232: data <= 8'h00;
            16'd4233: data <= 8'hF8;
            16'd4234: data <= 8'h00;
            16'd4235: data <= 8'hF8;
            16'd4236: data <= 8'h00;
            16'd4237: data <= 8'hF8;
            16'd4238: data <= 8'h00;
            16'd4239: data <= 8'hF8;
            16'd4240: data <= 8'hFF;
            16'd4241: data <= 8'hFF;
            16'd4242: data <= 8'h00;
            16'd4243: data <= 8'hF8;
            16'd4244: data <= 8'h00;
            16'd4245: data <= 8'hF8;
            16'd4246: data <= 8'h00;
            16'd4247: data <= 8'hF8;
            16'd4248: data <= 8'h00;
            16'd4249: data <= 8'hF8;
            16'd4250: data <= 8'h00;
            16'd4251: data <= 8'hF8;
            16'd4252: data <= 8'h00;
            16'd4253: data <= 8'hF8;
            16'd4254: data <= 8'h00;
            16'd4255: data <= 8'hF8;
            16'd4256: data <= 8'h00;
            16'd4257: data <= 8'hF8;
            16'd4258: data <= 8'h00;
            16'd4259: data <= 8'hF8;
            16'd4260: data <= 8'h00;
            16'd4261: data <= 8'hF8;
            16'd4262: data <= 8'h00;
            16'd4263: data <= 8'hF8;
            16'd4264: data <= 8'h00;
            16'd4265: data <= 8'hF8;
            16'd4266: data <= 8'h00;
            16'd4267: data <= 8'hF8;
            16'd4268: data <= 8'h00;
            16'd4269: data <= 8'hF8;
            16'd4270: data <= 8'h00;
            16'd4271: data <= 8'hF8;
            16'd4272: data <= 8'h00;
            16'd4273: data <= 8'hF8;
            16'd4274: data <= 8'h00;
            16'd4275: data <= 8'hF8;
            16'd4276: data <= 8'h00;
            16'd4277: data <= 8'hF8;
            16'd4278: data <= 8'h00;
            16'd4279: data <= 8'hF8;
            16'd4280: data <= 8'hFF;
            16'd4281: data <= 8'hFF;
            16'd4282: data <= 8'h00;
            16'd4283: data <= 8'hF8;
            16'd4284: data <= 8'h00;
            16'd4285: data <= 8'hF8;
            16'd4286: data <= 8'h00;
            16'd4287: data <= 8'hF8;
            16'd4288: data <= 8'h00;
            16'd4289: data <= 8'hF8;
            16'd4290: data <= 8'h00;
            16'd4291: data <= 8'hF8;
            16'd4292: data <= 8'h00;
            16'd4293: data <= 8'hF8;
            16'd4294: data <= 8'h00;
            16'd4295: data <= 8'hF8;
            16'd4296: data <= 8'h00;
            16'd4297: data <= 8'hF8;
            16'd4298: data <= 8'h00;
            16'd4299: data <= 8'hF8;
            16'd4300: data <= 8'h00;
            16'd4301: data <= 8'hF8;
            16'd4302: data <= 8'h00;
            16'd4303: data <= 8'hF8;
            16'd4304: data <= 8'h00;
            16'd4305: data <= 8'hF8;
            16'd4306: data <= 8'h00;
            16'd4307: data <= 8'hF8;
            16'd4308: data <= 8'h00;
            16'd4309: data <= 8'hF8;
            16'd4310: data <= 8'h00;
            16'd4311: data <= 8'hF8;
            16'd4312: data <= 8'h00;
            16'd4313: data <= 8'hF8;
            16'd4314: data <= 8'h00;
            16'd4315: data <= 8'hF8;
            16'd4316: data <= 8'h00;
            16'd4317: data <= 8'hF8;
            16'd4318: data <= 8'h00;
            16'd4319: data <= 8'hF8;
            16'd4320: data <= 8'hFF;
            16'd4321: data <= 8'hFF;
            16'd4322: data <= 8'h00;
            16'd4323: data <= 8'hF8;
            16'd4324: data <= 8'h00;
            16'd4325: data <= 8'hF8;
            16'd4326: data <= 8'h00;
            16'd4327: data <= 8'hF8;
            16'd4328: data <= 8'h00;
            16'd4329: data <= 8'hF8;
            16'd4330: data <= 8'h00;
            16'd4331: data <= 8'hF8;
            16'd4332: data <= 8'h00;
            16'd4333: data <= 8'hF8;
            16'd4334: data <= 8'h00;
            16'd4335: data <= 8'hF8;
            16'd4336: data <= 8'h00;
            16'd4337: data <= 8'hF8;
            16'd4338: data <= 8'h00;
            16'd4339: data <= 8'hF8;
            16'd4340: data <= 8'h00;
            16'd4341: data <= 8'hF8;
            16'd4342: data <= 8'h00;
            16'd4343: data <= 8'hF8;
            16'd4344: data <= 8'h00;
            16'd4345: data <= 8'hF8;
            16'd4346: data <= 8'h00;
            16'd4347: data <= 8'hF8;
            16'd4348: data <= 8'h00;
            16'd4349: data <= 8'hF8;
            16'd4350: data <= 8'h00;
            16'd4351: data <= 8'hF8;
            16'd4352: data <= 8'h00;
            16'd4353: data <= 8'hF8;
            16'd4354: data <= 8'h00;
            16'd4355: data <= 8'hF8;
            16'd4356: data <= 8'h00;
            16'd4357: data <= 8'hF8;
            16'd4358: data <= 8'h00;
            16'd4359: data <= 8'hF8;
            16'd4360: data <= 8'hFF;
            16'd4361: data <= 8'hFF;
            16'd4362: data <= 8'h00;
            16'd4363: data <= 8'hF8;
            16'd4364: data <= 8'h00;
            16'd4365: data <= 8'hF8;
            16'd4366: data <= 8'h00;
            16'd4367: data <= 8'hF8;
            16'd4368: data <= 8'h00;
            16'd4369: data <= 8'hF8;
            16'd4370: data <= 8'h00;
            16'd4371: data <= 8'hF8;
            16'd4372: data <= 8'h00;
            16'd4373: data <= 8'hF8;
            16'd4374: data <= 8'h00;
            16'd4375: data <= 8'hF8;
            16'd4376: data <= 8'h00;
            16'd4377: data <= 8'hF8;
            16'd4378: data <= 8'h00;
            16'd4379: data <= 8'hF8;
            16'd4380: data <= 8'h00;
            16'd4381: data <= 8'hF8;
            16'd4382: data <= 8'h00;
            16'd4383: data <= 8'hF8;
            16'd4384: data <= 8'h00;
            16'd4385: data <= 8'hF8;
            16'd4386: data <= 8'h00;
            16'd4387: data <= 8'hF8;
            16'd4388: data <= 8'h00;
            16'd4389: data <= 8'hF8;
            16'd4390: data <= 8'h00;
            16'd4391: data <= 8'hF8;
            16'd4392: data <= 8'h00;
            16'd4393: data <= 8'hF8;
            16'd4394: data <= 8'h00;
            16'd4395: data <= 8'hF8;
            16'd4396: data <= 8'h00;
            16'd4397: data <= 8'hF8;
            16'd4398: data <= 8'h00;
            16'd4399: data <= 8'hF8;
            16'd4400: data <= 8'hFF;
            16'd4401: data <= 8'hFF;
            16'd4402: data <= 8'h00;
            16'd4403: data <= 8'hF8;
            16'd4404: data <= 8'h00;
            16'd4405: data <= 8'hF8;
            16'd4406: data <= 8'h00;
            16'd4407: data <= 8'hF8;
            16'd4408: data <= 8'h00;
            16'd4409: data <= 8'hF8;
            16'd4410: data <= 8'h00;
            16'd4411: data <= 8'hF8;
            16'd4412: data <= 8'h00;
            16'd4413: data <= 8'hF8;
            16'd4414: data <= 8'h00;
            16'd4415: data <= 8'hF8;
            16'd4416: data <= 8'h00;
            16'd4417: data <= 8'hF8;
            16'd4418: data <= 8'h00;
            16'd4419: data <= 8'hF8;
            16'd4420: data <= 8'h00;
            16'd4421: data <= 8'hF8;
            16'd4422: data <= 8'h00;
            16'd4423: data <= 8'hF8;
            16'd4424: data <= 8'h00;
            16'd4425: data <= 8'hF8;
            16'd4426: data <= 8'h00;
            16'd4427: data <= 8'hF8;
            16'd4428: data <= 8'h00;
            16'd4429: data <= 8'hF8;
            16'd4430: data <= 8'h00;
            16'd4431: data <= 8'hF8;
            16'd4432: data <= 8'h00;
            16'd4433: data <= 8'hF8;
            16'd4434: data <= 8'h00;
            16'd4435: data <= 8'hF8;
            16'd4436: data <= 8'h00;
            16'd4437: data <= 8'hF8;
            16'd4438: data <= 8'h00;
            16'd4439: data <= 8'hF8;
            16'd4440: data <= 8'hFF;
            16'd4441: data <= 8'hFF;
            16'd4442: data <= 8'h00;
            16'd4443: data <= 8'hF8;
            16'd4444: data <= 8'h00;
            16'd4445: data <= 8'hF8;
            16'd4446: data <= 8'h00;
            16'd4447: data <= 8'hF8;
            16'd4448: data <= 8'h00;
            16'd4449: data <= 8'hF8;
            16'd4450: data <= 8'h00;
            16'd4451: data <= 8'hF8;
            16'd4452: data <= 8'h00;
            16'd4453: data <= 8'hF8;
            16'd4454: data <= 8'h00;
            16'd4455: data <= 8'hF8;
            16'd4456: data <= 8'h00;
            16'd4457: data <= 8'hF8;
            16'd4458: data <= 8'h00;
            16'd4459: data <= 8'hF8;
            16'd4460: data <= 8'h00;
            16'd4461: data <= 8'hF8;
            16'd4462: data <= 8'h00;
            16'd4463: data <= 8'hF8;
            16'd4464: data <= 8'h00;
            16'd4465: data <= 8'hF8;
            16'd4466: data <= 8'h00;
            16'd4467: data <= 8'hF8;
            16'd4468: data <= 8'h00;
            16'd4469: data <= 8'hF8;
            16'd4470: data <= 8'h00;
            16'd4471: data <= 8'hF8;
            16'd4472: data <= 8'h00;
            16'd4473: data <= 8'hF8;
            16'd4474: data <= 8'h00;
            16'd4475: data <= 8'hF8;
            16'd4476: data <= 8'h00;
            16'd4477: data <= 8'hF8;
            16'd4478: data <= 8'h00;
            16'd4479: data <= 8'hF8;
            16'd4480: data <= 8'hFF;
            16'd4481: data <= 8'hFF;
            16'd4482: data <= 8'h00;
            16'd4483: data <= 8'hF8;
            16'd4484: data <= 8'h00;
            16'd4485: data <= 8'hF8;
            16'd4486: data <= 8'h00;
            16'd4487: data <= 8'hF8;
            16'd4488: data <= 8'h00;
            16'd4489: data <= 8'hF8;
            16'd4490: data <= 8'h00;
            16'd4491: data <= 8'hF8;
            16'd4492: data <= 8'h00;
            16'd4493: data <= 8'hF8;
            16'd4494: data <= 8'h00;
            16'd4495: data <= 8'hF8;
            16'd4496: data <= 8'h00;
            16'd4497: data <= 8'hF8;
            16'd4498: data <= 8'h00;
            16'd4499: data <= 8'hF8;
            16'd4500: data <= 8'h00;
            16'd4501: data <= 8'hF8;
            16'd4502: data <= 8'h00;
            16'd4503: data <= 8'hF8;
            16'd4504: data <= 8'h00;
            16'd4505: data <= 8'hF8;
            16'd4506: data <= 8'h00;
            16'd4507: data <= 8'hF8;
            16'd4508: data <= 8'h00;
            16'd4509: data <= 8'hF8;
            16'd4510: data <= 8'h00;
            16'd4511: data <= 8'hF8;
            16'd4512: data <= 8'h00;
            16'd4513: data <= 8'hF8;
            16'd4514: data <= 8'h00;
            16'd4515: data <= 8'hF8;
            16'd4516: data <= 8'h00;
            16'd4517: data <= 8'hF8;
            16'd4518: data <= 8'h00;
            16'd4519: data <= 8'hF8;
            16'd4520: data <= 8'hFF;
            16'd4521: data <= 8'hFF;
            16'd4522: data <= 8'h00;
            16'd4523: data <= 8'hF8;
            16'd4524: data <= 8'h00;
            16'd4525: data <= 8'hF8;
            16'd4526: data <= 8'h00;
            16'd4527: data <= 8'hF8;
            16'd4528: data <= 8'h00;
            16'd4529: data <= 8'hF8;
            16'd4530: data <= 8'h00;
            16'd4531: data <= 8'hF8;
            16'd4532: data <= 8'h00;
            16'd4533: data <= 8'hF8;
            16'd4534: data <= 8'h00;
            16'd4535: data <= 8'hF8;
            16'd4536: data <= 8'h00;
            16'd4537: data <= 8'hF8;
            16'd4538: data <= 8'h00;
            16'd4539: data <= 8'hF8;
            16'd4540: data <= 8'h00;
            16'd4541: data <= 8'hF8;
            16'd4542: data <= 8'h00;
            16'd4543: data <= 8'hF8;
            16'd4544: data <= 8'h00;
            16'd4545: data <= 8'hF8;
            16'd4546: data <= 8'h00;
            16'd4547: data <= 8'hF8;
            16'd4548: data <= 8'h00;
            16'd4549: data <= 8'hF8;
            16'd4550: data <= 8'h00;
            16'd4551: data <= 8'hF8;
            16'd4552: data <= 8'h00;
            16'd4553: data <= 8'hF8;
            16'd4554: data <= 8'h00;
            16'd4555: data <= 8'hF8;
            16'd4556: data <= 8'h00;
            16'd4557: data <= 8'hF8;
            16'd4558: data <= 8'h00;
            16'd4559: data <= 8'hF8;
            16'd4560: data <= 8'hFF;
            16'd4561: data <= 8'hFF;
            16'd4562: data <= 8'h00;
            16'd4563: data <= 8'hF8;
            16'd4564: data <= 8'h00;
            16'd4565: data <= 8'hF8;
            16'd4566: data <= 8'h00;
            16'd4567: data <= 8'hF8;
            16'd4568: data <= 8'h00;
            16'd4569: data <= 8'hF8;
            16'd4570: data <= 8'h00;
            16'd4571: data <= 8'hF8;
            16'd4572: data <= 8'h00;
            16'd4573: data <= 8'hF8;
            16'd4574: data <= 8'h00;
            16'd4575: data <= 8'hF8;
            16'd4576: data <= 8'h00;
            16'd4577: data <= 8'hF8;
            16'd4578: data <= 8'h00;
            16'd4579: data <= 8'hF8;
            16'd4580: data <= 8'h00;
            16'd4581: data <= 8'hF8;
            16'd4582: data <= 8'h00;
            16'd4583: data <= 8'hF8;
            16'd4584: data <= 8'h00;
            16'd4585: data <= 8'hF8;
            16'd4586: data <= 8'h00;
            16'd4587: data <= 8'hF8;
            16'd4588: data <= 8'h00;
            16'd4589: data <= 8'hF8;
            16'd4590: data <= 8'h00;
            16'd4591: data <= 8'hF8;
            16'd4592: data <= 8'h00;
            16'd4593: data <= 8'hF8;
            16'd4594: data <= 8'h00;
            16'd4595: data <= 8'hF8;
            16'd4596: data <= 8'h00;
            16'd4597: data <= 8'hF8;
            16'd4598: data <= 8'h00;
            16'd4599: data <= 8'hF8;
            16'd4600: data <= 8'hFF;
            16'd4601: data <= 8'hFF;
            16'd4602: data <= 8'h00;
            16'd4603: data <= 8'hF8;
            16'd4604: data <= 8'h00;
            16'd4605: data <= 8'hF8;
            16'd4606: data <= 8'h00;
            16'd4607: data <= 8'hF8;
            16'd4608: data <= 8'h00;
            16'd4609: data <= 8'hF8;
            16'd4610: data <= 8'h00;
            16'd4611: data <= 8'hF8;
            16'd4612: data <= 8'h00;
            16'd4613: data <= 8'hF8;
            16'd4614: data <= 8'h00;
            16'd4615: data <= 8'hF8;
            16'd4616: data <= 8'h00;
            16'd4617: data <= 8'hF8;
            16'd4618: data <= 8'h00;
            16'd4619: data <= 8'hF8;
            16'd4620: data <= 8'h00;
            16'd4621: data <= 8'hF8;
            16'd4622: data <= 8'h00;
            16'd4623: data <= 8'hF8;
            16'd4624: data <= 8'h00;
            16'd4625: data <= 8'hF8;
            16'd4626: data <= 8'h00;
            16'd4627: data <= 8'hF8;
            16'd4628: data <= 8'h00;
            16'd4629: data <= 8'hF8;
            16'd4630: data <= 8'h00;
            16'd4631: data <= 8'hF8;
            16'd4632: data <= 8'h00;
            16'd4633: data <= 8'hF8;
            16'd4634: data <= 8'h00;
            16'd4635: data <= 8'hF8;
            16'd4636: data <= 8'h00;
            16'd4637: data <= 8'hF8;
            16'd4638: data <= 8'h00;
            16'd4639: data <= 8'hF8;
            16'd4640: data <= 8'hFF;
            16'd4641: data <= 8'hFF;
            16'd4642: data <= 8'h00;
            16'd4643: data <= 8'hF8;
            16'd4644: data <= 8'h00;
            16'd4645: data <= 8'hF8;
            16'd4646: data <= 8'h00;
            16'd4647: data <= 8'hF8;
            16'd4648: data <= 8'h00;
            16'd4649: data <= 8'hF8;
            16'd4650: data <= 8'h00;
            16'd4651: data <= 8'hF8;
            16'd4652: data <= 8'h00;
            16'd4653: data <= 8'hF8;
            16'd4654: data <= 8'h00;
            16'd4655: data <= 8'hF8;
            16'd4656: data <= 8'h00;
            16'd4657: data <= 8'hF8;
            16'd4658: data <= 8'h00;
            16'd4659: data <= 8'hF8;
            16'd4660: data <= 8'h00;
            16'd4661: data <= 8'hF8;
            16'd4662: data <= 8'h00;
            16'd4663: data <= 8'hF8;
            16'd4664: data <= 8'h00;
            16'd4665: data <= 8'hF8;
            16'd4666: data <= 8'h00;
            16'd4667: data <= 8'hF8;
            16'd4668: data <= 8'h00;
            16'd4669: data <= 8'hF8;
            16'd4670: data <= 8'h00;
            16'd4671: data <= 8'hF8;
            16'd4672: data <= 8'h00;
            16'd4673: data <= 8'hF8;
            16'd4674: data <= 8'h00;
            16'd4675: data <= 8'hF8;
            16'd4676: data <= 8'h00;
            16'd4677: data <= 8'hF8;
            16'd4678: data <= 8'h00;
            16'd4679: data <= 8'hF8;
            16'd4680: data <= 8'hFF;
            16'd4681: data <= 8'hFF;
            16'd4682: data <= 8'h00;
            16'd4683: data <= 8'hF8;
            16'd4684: data <= 8'h00;
            16'd4685: data <= 8'hF8;
            16'd4686: data <= 8'h00;
            16'd4687: data <= 8'hF8;
            16'd4688: data <= 8'h00;
            16'd4689: data <= 8'hF8;
            16'd4690: data <= 8'h00;
            16'd4691: data <= 8'hF8;
            16'd4692: data <= 8'h00;
            16'd4693: data <= 8'hF8;
            16'd4694: data <= 8'h00;
            16'd4695: data <= 8'hF8;
            16'd4696: data <= 8'h00;
            16'd4697: data <= 8'hF8;
            16'd4698: data <= 8'h00;
            16'd4699: data <= 8'hF8;
            16'd4700: data <= 8'h00;
            16'd4701: data <= 8'hF8;
            16'd4702: data <= 8'h00;
            16'd4703: data <= 8'hF8;
            16'd4704: data <= 8'h00;
            16'd4705: data <= 8'hF8;
            16'd4706: data <= 8'h00;
            16'd4707: data <= 8'hF8;
            16'd4708: data <= 8'h00;
            16'd4709: data <= 8'hF8;
            16'd4710: data <= 8'h00;
            16'd4711: data <= 8'hF8;
            16'd4712: data <= 8'h00;
            16'd4713: data <= 8'hF8;
            16'd4714: data <= 8'h00;
            16'd4715: data <= 8'hF8;
            16'd4716: data <= 8'h00;
            16'd4717: data <= 8'hF8;
            16'd4718: data <= 8'h00;
            16'd4719: data <= 8'hF8;
            16'd4720: data <= 8'hFF;
            16'd4721: data <= 8'hFF;
            16'd4722: data <= 8'h00;
            16'd4723: data <= 8'hF8;
            16'd4724: data <= 8'h00;
            16'd4725: data <= 8'hF8;
            16'd4726: data <= 8'h00;
            16'd4727: data <= 8'hF8;
            16'd4728: data <= 8'h00;
            16'd4729: data <= 8'hF8;
            16'd4730: data <= 8'h00;
            16'd4731: data <= 8'hF8;
            16'd4732: data <= 8'h00;
            16'd4733: data <= 8'hF8;
            16'd4734: data <= 8'h00;
            16'd4735: data <= 8'hF8;
            16'd4736: data <= 8'h00;
            16'd4737: data <= 8'hF8;
            16'd4738: data <= 8'h00;
            16'd4739: data <= 8'hF8;
            16'd4740: data <= 8'h00;
            16'd4741: data <= 8'hF8;
            16'd4742: data <= 8'h00;
            16'd4743: data <= 8'hF8;
            16'd4744: data <= 8'h00;
            16'd4745: data <= 8'hF8;
            16'd4746: data <= 8'h00;
            16'd4747: data <= 8'hF8;
            16'd4748: data <= 8'h00;
            16'd4749: data <= 8'hF8;
            16'd4750: data <= 8'h00;
            16'd4751: data <= 8'hF8;
            16'd4752: data <= 8'h00;
            16'd4753: data <= 8'hF8;
            16'd4754: data <= 8'h00;
            16'd4755: data <= 8'hF8;
            16'd4756: data <= 8'h00;
            16'd4757: data <= 8'hF8;
            16'd4758: data <= 8'h00;
            16'd4759: data <= 8'hF8;
            16'd4760: data <= 8'hFF;
            16'd4761: data <= 8'hFF;
            16'd4762: data <= 8'h00;
            16'd4763: data <= 8'hF8;
            16'd4764: data <= 8'h00;
            16'd4765: data <= 8'hF8;
            16'd4766: data <= 8'h00;
            16'd4767: data <= 8'hF8;
            16'd4768: data <= 8'h00;
            16'd4769: data <= 8'hF8;
            16'd4770: data <= 8'h00;
            16'd4771: data <= 8'hF8;
            16'd4772: data <= 8'h00;
            16'd4773: data <= 8'hF8;
            16'd4774: data <= 8'h00;
            16'd4775: data <= 8'hF8;
            16'd4776: data <= 8'h00;
            16'd4777: data <= 8'hF8;
            16'd4778: data <= 8'h00;
            16'd4779: data <= 8'hF8;
            16'd4780: data <= 8'h00;
            16'd4781: data <= 8'hF8;
            16'd4782: data <= 8'h00;
            16'd4783: data <= 8'hF8;
            16'd4784: data <= 8'h00;
            16'd4785: data <= 8'hF8;
            16'd4786: data <= 8'h00;
            16'd4787: data <= 8'hF8;
            16'd4788: data <= 8'h00;
            16'd4789: data <= 8'hF8;
            16'd4790: data <= 8'h00;
            16'd4791: data <= 8'hF8;
            16'd4792: data <= 8'h00;
            16'd4793: data <= 8'hF8;
            16'd4794: data <= 8'h00;
            16'd4795: data <= 8'hF8;
            16'd4796: data <= 8'h00;
            16'd4797: data <= 8'hF8;
            16'd4798: data <= 8'h00;
            16'd4799: data <= 8'hF8;
            16'd4800: data <= 8'hFF;
            16'd4801: data <= 8'hFF;
            16'd4802: data <= 8'hFF;
            16'd4803: data <= 8'hFF;
            16'd4804: data <= 8'hFF;
            16'd4805: data <= 8'hFF;
            16'd4806: data <= 8'hFF;
            16'd4807: data <= 8'hFF;
            16'd4808: data <= 8'hFF;
            16'd4809: data <= 8'hFF;
            16'd4810: data <= 8'hFF;
            16'd4811: data <= 8'hFF;
            16'd4812: data <= 8'hFF;
            16'd4813: data <= 8'hFF;
            16'd4814: data <= 8'hFF;
            16'd4815: data <= 8'hFF;
            16'd4816: data <= 8'hFF;
            16'd4817: data <= 8'hFF;
            16'd4818: data <= 8'hFF;
            16'd4819: data <= 8'hFF;
            16'd4820: data <= 8'hFF;
            16'd4821: data <= 8'hFF;
            16'd4822: data <= 8'hFF;
            16'd4823: data <= 8'hFF;
            16'd4824: data <= 8'hFF;
            16'd4825: data <= 8'hFF;
            16'd4826: data <= 8'hFF;
            16'd4827: data <= 8'hFF;
            16'd4828: data <= 8'hFF;
            16'd4829: data <= 8'hFF;
            16'd4830: data <= 8'hFF;
            16'd4831: data <= 8'hFF;
            16'd4832: data <= 8'hFF;
            16'd4833: data <= 8'hFF;
            16'd4834: data <= 8'hFF;
            16'd4835: data <= 8'hFF;
            16'd4836: data <= 8'hFF;
            16'd4837: data <= 8'hFF;
            16'd4838: data <= 8'hFF;
            16'd4839: data <= 8'hFF;
            16'd4840: data <= 8'hFF;
            16'd4841: data <= 8'hFF;
            16'd4842: data <= 8'hFF;
            16'd4843: data <= 8'hFF;
            16'd4844: data <= 8'hFF;
            16'd4845: data <= 8'hFF;
            16'd4846: data <= 8'hFF;
            16'd4847: data <= 8'hFF;
            16'd4848: data <= 8'hFF;
            16'd4849: data <= 8'hFF;
            16'd4850: data <= 8'hFF;
            16'd4851: data <= 8'hFF;
            16'd4852: data <= 8'hFF;
            16'd4853: data <= 8'hFF;
            16'd4854: data <= 8'hFF;
            16'd4855: data <= 8'hFF;
            16'd4856: data <= 8'hFF;
            16'd4857: data <= 8'hFF;
            16'd4858: data <= 8'hFF;
            16'd4859: data <= 8'hFF;
            16'd4860: data <= 8'hFF;
            16'd4861: data <= 8'hFF;
            16'd4862: data <= 8'hFF;
            16'd4863: data <= 8'hFF;
            16'd4864: data <= 8'hFF;
            16'd4865: data <= 8'hFF;
            16'd4866: data <= 8'hFF;
            16'd4867: data <= 8'hFF;
            16'd4868: data <= 8'hFF;
            16'd4869: data <= 8'hFF;
            16'd4870: data <= 8'hFF;
            16'd4871: data <= 8'hFF;
            16'd4872: data <= 8'hFF;
            16'd4873: data <= 8'hFF;
            16'd4874: data <= 8'hFF;
            16'd4875: data <= 8'hFF;
            16'd4876: data <= 8'hFF;
            16'd4877: data <= 8'hFF;
            16'd4878: data <= 8'hFF;
            16'd4879: data <= 8'hFF;
            16'd4880: data <= 8'hFF;
            16'd4881: data <= 8'hFF;
            16'd4882: data <= 8'hFF;
            16'd4883: data <= 8'hFF;
            16'd4884: data <= 8'hFF;
            16'd4885: data <= 8'hFF;
            16'd4886: data <= 8'hFF;
            16'd4887: data <= 8'hFF;
            16'd4888: data <= 8'hFF;
            16'd4889: data <= 8'hFF;
            16'd4890: data <= 8'hFF;
            16'd4891: data <= 8'hFF;
            16'd4892: data <= 8'hFF;
            16'd4893: data <= 8'hFF;
            16'd4894: data <= 8'hFF;
            16'd4895: data <= 8'hFF;
            16'd4896: data <= 8'hFF;
            16'd4897: data <= 8'hFF;
            16'd4898: data <= 8'hFF;
            16'd4899: data <= 8'hFF;
            16'd4900: data <= 8'hFF;
            16'd4901: data <= 8'hFF;
            16'd4902: data <= 8'hFF;
            16'd4903: data <= 8'hFF;
            16'd4904: data <= 8'hFF;
            16'd4905: data <= 8'hFF;
            16'd4906: data <= 8'hFF;
            16'd4907: data <= 8'hFF;
            16'd4908: data <= 8'hFF;
            16'd4909: data <= 8'hFF;
            16'd4910: data <= 8'hFF;
            16'd4911: data <= 8'hFF;
            16'd4912: data <= 8'hFF;
            16'd4913: data <= 8'hFF;
            16'd4914: data <= 8'hFF;
            16'd4915: data <= 8'hFF;
            16'd4916: data <= 8'hFF;
            16'd4917: data <= 8'hFF;
            16'd4918: data <= 8'hFF;
            16'd4919: data <= 8'hFF;
            16'd4920: data <= 8'hFF;
            16'd4921: data <= 8'hFF;
            16'd4922: data <= 8'hFF;
            16'd4923: data <= 8'hFF;
            16'd4924: data <= 8'hFF;
            16'd4925: data <= 8'hFF;
            16'd4926: data <= 8'hFF;
            16'd4927: data <= 8'hFF;
            16'd4928: data <= 8'hFF;
            16'd4929: data <= 8'hFF;
            16'd4930: data <= 8'hFF;
            16'd4931: data <= 8'hFF;
            16'd4932: data <= 8'hFF;
            16'd4933: data <= 8'hFF;
            16'd4934: data <= 8'hFF;
            16'd4935: data <= 8'hFF;
            16'd4936: data <= 8'hFF;
            16'd4937: data <= 8'hFF;
            16'd4938: data <= 8'hFF;
            16'd4939: data <= 8'hFF;
            16'd4940: data <= 8'hFF;
            16'd4941: data <= 8'hFF;
            16'd4942: data <= 8'hFF;
            16'd4943: data <= 8'hFF;
            16'd4944: data <= 8'hFF;
            16'd4945: data <= 8'hFF;
            16'd4946: data <= 8'hFF;
            16'd4947: data <= 8'hFF;
            16'd4948: data <= 8'hFF;
            16'd4949: data <= 8'hFF;
            16'd4950: data <= 8'hFF;
            16'd4951: data <= 8'hFF;
            16'd4952: data <= 8'hFF;
            16'd4953: data <= 8'hFF;
            16'd4954: data <= 8'hFF;
            16'd4955: data <= 8'hFF;
            16'd4956: data <= 8'hFF;
            16'd4957: data <= 8'hFF;
            16'd4958: data <= 8'hFF;
            16'd4959: data <= 8'hFF;
            16'd4960: data <= 8'hFF;
            16'd4961: data <= 8'hFF;
            16'd4962: data <= 8'hFF;
            16'd4963: data <= 8'hFF;
            16'd4964: data <= 8'hFF;
            16'd4965: data <= 8'hFF;
            16'd4966: data <= 8'hFF;
            16'd4967: data <= 8'hFF;
            16'd4968: data <= 8'hFF;
            16'd4969: data <= 8'hFF;
            16'd4970: data <= 8'hFF;
            16'd4971: data <= 8'hFF;
            16'd4972: data <= 8'hFF;
            16'd4973: data <= 8'hFF;
            16'd4974: data <= 8'hFF;
            16'd4975: data <= 8'hFF;
            16'd4976: data <= 8'hFF;
            16'd4977: data <= 8'hFF;
            16'd4978: data <= 8'hFF;
            16'd4979: data <= 8'hFF;
            16'd4980: data <= 8'hFF;
            16'd4981: data <= 8'hFF;
            16'd4982: data <= 8'hFF;
            16'd4983: data <= 8'hFF;
            16'd4984: data <= 8'hFF;
            16'd4985: data <= 8'hFF;
            16'd4986: data <= 8'hFF;
            16'd4987: data <= 8'hFF;
            16'd4988: data <= 8'hFF;
            16'd4989: data <= 8'hFF;
            16'd4990: data <= 8'hFF;
            16'd4991: data <= 8'hFF;
            16'd4992: data <= 8'hFF;
            16'd4993: data <= 8'hFF;
            16'd4994: data <= 8'hFF;
            16'd4995: data <= 8'hFF;
            16'd4996: data <= 8'hFF;
            16'd4997: data <= 8'hFF;
            16'd4998: data <= 8'hFF;
            16'd4999: data <= 8'hFF;
            16'd5000: data <= 8'hFF;
            16'd5001: data <= 8'hFF;
            16'd5002: data <= 8'hFF;
            16'd5003: data <= 8'hFF;
            16'd5004: data <= 8'hFF;
            16'd5005: data <= 8'hFF;
            16'd5006: data <= 8'hFF;
            16'd5007: data <= 8'hFF;
            16'd5008: data <= 8'hFF;
            16'd5009: data <= 8'hFF;
            16'd5010: data <= 8'hFF;
            16'd5011: data <= 8'hFF;
            16'd5012: data <= 8'hFF;
            16'd5013: data <= 8'hFF;
            16'd5014: data <= 8'hFF;
            16'd5015: data <= 8'hFF;
            16'd5016: data <= 8'hFF;
            16'd5017: data <= 8'hFF;
            16'd5018: data <= 8'hFF;
            16'd5019: data <= 8'hFF;
            16'd5020: data <= 8'hFF;
            16'd5021: data <= 8'hFF;
            16'd5022: data <= 8'hFF;
            16'd5023: data <= 8'hFF;
            16'd5024: data <= 8'hFF;
            16'd5025: data <= 8'hFF;
            16'd5026: data <= 8'hFF;
            16'd5027: data <= 8'hFF;
            16'd5028: data <= 8'hFF;
            16'd5029: data <= 8'hFF;
            16'd5030: data <= 8'hFF;
            16'd5031: data <= 8'hFF;
            16'd5032: data <= 8'hFF;
            16'd5033: data <= 8'hFF;
            16'd5034: data <= 8'hFF;
            16'd5035: data <= 8'hFF;
            16'd5036: data <= 8'hFF;
            16'd5037: data <= 8'hFF;
            16'd5038: data <= 8'hFF;
            16'd5039: data <= 8'hFF;
            16'd5040: data <= 8'hFF;
            16'd5041: data <= 8'hFF;
            16'd5042: data <= 8'h00;
            16'd5043: data <= 8'hF8;
            16'd5044: data <= 8'h00;
            16'd5045: data <= 8'hF8;
            16'd5046: data <= 8'h00;
            16'd5047: data <= 8'hF8;
            16'd5048: data <= 8'h00;
            16'd5049: data <= 8'hF8;
            16'd5050: data <= 8'h00;
            16'd5051: data <= 8'hF8;
            16'd5052: data <= 8'h00;
            16'd5053: data <= 8'hF8;
            16'd5054: data <= 8'h00;
            16'd5055: data <= 8'hF8;
            16'd5056: data <= 8'h00;
            16'd5057: data <= 8'hF8;
            16'd5058: data <= 8'h00;
            16'd5059: data <= 8'hF8;
            16'd5060: data <= 8'h00;
            16'd5061: data <= 8'hF8;
            16'd5062: data <= 8'h00;
            16'd5063: data <= 8'hF8;
            16'd5064: data <= 8'h00;
            16'd5065: data <= 8'hF8;
            16'd5066: data <= 8'h00;
            16'd5067: data <= 8'hF8;
            16'd5068: data <= 8'h00;
            16'd5069: data <= 8'hF8;
            16'd5070: data <= 8'h00;
            16'd5071: data <= 8'hF8;
            16'd5072: data <= 8'h00;
            16'd5073: data <= 8'hF8;
            16'd5074: data <= 8'h00;
            16'd5075: data <= 8'hF8;
            16'd5076: data <= 8'h00;
            16'd5077: data <= 8'hF8;
            16'd5078: data <= 8'h00;
            16'd5079: data <= 8'hF8;
            16'd5080: data <= 8'hFF;
            16'd5081: data <= 8'hFF;
            16'd5082: data <= 8'h00;
            16'd5083: data <= 8'hF8;
            16'd5084: data <= 8'h00;
            16'd5085: data <= 8'hF8;
            16'd5086: data <= 8'h00;
            16'd5087: data <= 8'hF8;
            16'd5088: data <= 8'h00;
            16'd5089: data <= 8'hF8;
            16'd5090: data <= 8'h00;
            16'd5091: data <= 8'hF8;
            16'd5092: data <= 8'h00;
            16'd5093: data <= 8'hF8;
            16'd5094: data <= 8'h00;
            16'd5095: data <= 8'hF8;
            16'd5096: data <= 8'h00;
            16'd5097: data <= 8'hF8;
            16'd5098: data <= 8'h00;
            16'd5099: data <= 8'hF8;
            16'd5100: data <= 8'h00;
            16'd5101: data <= 8'hF8;
            16'd5102: data <= 8'h00;
            16'd5103: data <= 8'hF8;
            16'd5104: data <= 8'h00;
            16'd5105: data <= 8'hF8;
            16'd5106: data <= 8'h00;
            16'd5107: data <= 8'hF8;
            16'd5108: data <= 8'h00;
            16'd5109: data <= 8'hF8;
            16'd5110: data <= 8'h00;
            16'd5111: data <= 8'hF8;
            16'd5112: data <= 8'h00;
            16'd5113: data <= 8'hF8;
            16'd5114: data <= 8'h00;
            16'd5115: data <= 8'hF8;
            16'd5116: data <= 8'h00;
            16'd5117: data <= 8'hF8;
            16'd5118: data <= 8'h00;
            16'd5119: data <= 8'hF8;
            16'd5120: data <= 8'hFF;
            16'd5121: data <= 8'hFF;
            16'd5122: data <= 8'h00;
            16'd5123: data <= 8'hF8;
            16'd5124: data <= 8'h00;
            16'd5125: data <= 8'hF8;
            16'd5126: data <= 8'h00;
            16'd5127: data <= 8'hF8;
            16'd5128: data <= 8'h00;
            16'd5129: data <= 8'hF8;
            16'd5130: data <= 8'h00;
            16'd5131: data <= 8'hF8;
            16'd5132: data <= 8'h00;
            16'd5133: data <= 8'hF8;
            16'd5134: data <= 8'h00;
            16'd5135: data <= 8'hF8;
            16'd5136: data <= 8'h00;
            16'd5137: data <= 8'hF8;
            16'd5138: data <= 8'h00;
            16'd5139: data <= 8'hF8;
            16'd5140: data <= 8'h00;
            16'd5141: data <= 8'hF8;
            16'd5142: data <= 8'h00;
            16'd5143: data <= 8'hF8;
            16'd5144: data <= 8'h00;
            16'd5145: data <= 8'hF8;
            16'd5146: data <= 8'h00;
            16'd5147: data <= 8'hF8;
            16'd5148: data <= 8'h00;
            16'd5149: data <= 8'hF8;
            16'd5150: data <= 8'h00;
            16'd5151: data <= 8'hF8;
            16'd5152: data <= 8'h00;
            16'd5153: data <= 8'hF8;
            16'd5154: data <= 8'h00;
            16'd5155: data <= 8'hF8;
            16'd5156: data <= 8'h00;
            16'd5157: data <= 8'hF8;
            16'd5158: data <= 8'h00;
            16'd5159: data <= 8'hF8;
            16'd5160: data <= 8'hFF;
            16'd5161: data <= 8'hFF;
            16'd5162: data <= 8'h00;
            16'd5163: data <= 8'hF8;
            16'd5164: data <= 8'h00;
            16'd5165: data <= 8'hF8;
            16'd5166: data <= 8'h00;
            16'd5167: data <= 8'hF8;
            16'd5168: data <= 8'h00;
            16'd5169: data <= 8'hF8;
            16'd5170: data <= 8'h00;
            16'd5171: data <= 8'hF8;
            16'd5172: data <= 8'h00;
            16'd5173: data <= 8'hF8;
            16'd5174: data <= 8'h00;
            16'd5175: data <= 8'hF8;
            16'd5176: data <= 8'h00;
            16'd5177: data <= 8'hF8;
            16'd5178: data <= 8'h00;
            16'd5179: data <= 8'hF8;
            16'd5180: data <= 8'h00;
            16'd5181: data <= 8'hF8;
            16'd5182: data <= 8'h00;
            16'd5183: data <= 8'hF8;
            16'd5184: data <= 8'h00;
            16'd5185: data <= 8'hF8;
            16'd5186: data <= 8'h00;
            16'd5187: data <= 8'hF8;
            16'd5188: data <= 8'h00;
            16'd5189: data <= 8'hF8;
            16'd5190: data <= 8'h00;
            16'd5191: data <= 8'hF8;
            16'd5192: data <= 8'h00;
            16'd5193: data <= 8'hF8;
            16'd5194: data <= 8'h00;
            16'd5195: data <= 8'hF8;
            16'd5196: data <= 8'h00;
            16'd5197: data <= 8'hF8;
            16'd5198: data <= 8'h00;
            16'd5199: data <= 8'hF8;
            16'd5200: data <= 8'hFF;
            16'd5201: data <= 8'hFF;
            16'd5202: data <= 8'h00;
            16'd5203: data <= 8'hF8;
            16'd5204: data <= 8'h00;
            16'd5205: data <= 8'hF8;
            16'd5206: data <= 8'h00;
            16'd5207: data <= 8'hF8;
            16'd5208: data <= 8'h00;
            16'd5209: data <= 8'hF8;
            16'd5210: data <= 8'h00;
            16'd5211: data <= 8'hF8;
            16'd5212: data <= 8'h00;
            16'd5213: data <= 8'hF8;
            16'd5214: data <= 8'h00;
            16'd5215: data <= 8'hF8;
            16'd5216: data <= 8'h00;
            16'd5217: data <= 8'hF8;
            16'd5218: data <= 8'h00;
            16'd5219: data <= 8'hF8;
            16'd5220: data <= 8'h00;
            16'd5221: data <= 8'hF8;
            16'd5222: data <= 8'h00;
            16'd5223: data <= 8'hF8;
            16'd5224: data <= 8'h00;
            16'd5225: data <= 8'hF8;
            16'd5226: data <= 8'h00;
            16'd5227: data <= 8'hF8;
            16'd5228: data <= 8'h00;
            16'd5229: data <= 8'hF8;
            16'd5230: data <= 8'h00;
            16'd5231: data <= 8'hF8;
            16'd5232: data <= 8'h00;
            16'd5233: data <= 8'hF8;
            16'd5234: data <= 8'h00;
            16'd5235: data <= 8'hF8;
            16'd5236: data <= 8'h00;
            16'd5237: data <= 8'hF8;
            16'd5238: data <= 8'h00;
            16'd5239: data <= 8'hF8;
            16'd5240: data <= 8'hFF;
            16'd5241: data <= 8'hFF;
            16'd5242: data <= 8'h00;
            16'd5243: data <= 8'hF8;
            16'd5244: data <= 8'h00;
            16'd5245: data <= 8'hF8;
            16'd5246: data <= 8'h00;
            16'd5247: data <= 8'hF8;
            16'd5248: data <= 8'h00;
            16'd5249: data <= 8'hF8;
            16'd5250: data <= 8'h00;
            16'd5251: data <= 8'hF8;
            16'd5252: data <= 8'h00;
            16'd5253: data <= 8'hF8;
            16'd5254: data <= 8'h00;
            16'd5255: data <= 8'hF8;
            16'd5256: data <= 8'h00;
            16'd5257: data <= 8'hF8;
            16'd5258: data <= 8'h00;
            16'd5259: data <= 8'hF8;
            16'd5260: data <= 8'h00;
            16'd5261: data <= 8'hF8;
            16'd5262: data <= 8'h00;
            16'd5263: data <= 8'hF8;
            16'd5264: data <= 8'h00;
            16'd5265: data <= 8'hF8;
            16'd5266: data <= 8'h00;
            16'd5267: data <= 8'hF8;
            16'd5268: data <= 8'h00;
            16'd5269: data <= 8'hF8;
            16'd5270: data <= 8'h00;
            16'd5271: data <= 8'hF8;
            16'd5272: data <= 8'h00;
            16'd5273: data <= 8'hF8;
            16'd5274: data <= 8'h00;
            16'd5275: data <= 8'hF8;
            16'd5276: data <= 8'h00;
            16'd5277: data <= 8'hF8;
            16'd5278: data <= 8'h00;
            16'd5279: data <= 8'hF8;
            16'd5280: data <= 8'hFF;
            16'd5281: data <= 8'hFF;
            16'd5282: data <= 8'h00;
            16'd5283: data <= 8'hF8;
            16'd5284: data <= 8'h00;
            16'd5285: data <= 8'hF8;
            16'd5286: data <= 8'h00;
            16'd5287: data <= 8'hF8;
            16'd5288: data <= 8'h00;
            16'd5289: data <= 8'hF8;
            16'd5290: data <= 8'h00;
            16'd5291: data <= 8'hF8;
            16'd5292: data <= 8'h00;
            16'd5293: data <= 8'hF8;
            16'd5294: data <= 8'h00;
            16'd5295: data <= 8'hF8;
            16'd5296: data <= 8'h00;
            16'd5297: data <= 8'hF8;
            16'd5298: data <= 8'h00;
            16'd5299: data <= 8'hF8;
            16'd5300: data <= 8'h00;
            16'd5301: data <= 8'hF8;
            16'd5302: data <= 8'h00;
            16'd5303: data <= 8'hF8;
            16'd5304: data <= 8'h00;
            16'd5305: data <= 8'hF8;
            16'd5306: data <= 8'h00;
            16'd5307: data <= 8'hF8;
            16'd5308: data <= 8'h00;
            16'd5309: data <= 8'hF8;
            16'd5310: data <= 8'h00;
            16'd5311: data <= 8'hF8;
            16'd5312: data <= 8'h00;
            16'd5313: data <= 8'hF8;
            16'd5314: data <= 8'h00;
            16'd5315: data <= 8'hF8;
            16'd5316: data <= 8'h00;
            16'd5317: data <= 8'hF8;
            16'd5318: data <= 8'h00;
            16'd5319: data <= 8'hF8;
            16'd5320: data <= 8'hFF;
            16'd5321: data <= 8'hFF;
            16'd5322: data <= 8'h00;
            16'd5323: data <= 8'hF8;
            16'd5324: data <= 8'h00;
            16'd5325: data <= 8'hF8;
            16'd5326: data <= 8'h00;
            16'd5327: data <= 8'hF8;
            16'd5328: data <= 8'h00;
            16'd5329: data <= 8'hF8;
            16'd5330: data <= 8'h00;
            16'd5331: data <= 8'hF8;
            16'd5332: data <= 8'h00;
            16'd5333: data <= 8'hF8;
            16'd5334: data <= 8'h00;
            16'd5335: data <= 8'hF8;
            16'd5336: data <= 8'h00;
            16'd5337: data <= 8'hF8;
            16'd5338: data <= 8'h00;
            16'd5339: data <= 8'hF8;
            16'd5340: data <= 8'h00;
            16'd5341: data <= 8'hF8;
            16'd5342: data <= 8'h00;
            16'd5343: data <= 8'hF8;
            16'd5344: data <= 8'h00;
            16'd5345: data <= 8'hF8;
            16'd5346: data <= 8'h00;
            16'd5347: data <= 8'hF8;
            16'd5348: data <= 8'h00;
            16'd5349: data <= 8'hF8;
            16'd5350: data <= 8'h00;
            16'd5351: data <= 8'hF8;
            16'd5352: data <= 8'h00;
            16'd5353: data <= 8'hF8;
            16'd5354: data <= 8'h00;
            16'd5355: data <= 8'hF8;
            16'd5356: data <= 8'h00;
            16'd5357: data <= 8'hF8;
            16'd5358: data <= 8'h00;
            16'd5359: data <= 8'hF8;
            16'd5360: data <= 8'hFF;
            16'd5361: data <= 8'hFF;
            16'd5362: data <= 8'h00;
            16'd5363: data <= 8'hF8;
            16'd5364: data <= 8'h00;
            16'd5365: data <= 8'hF8;
            16'd5366: data <= 8'h00;
            16'd5367: data <= 8'hF8;
            16'd5368: data <= 8'h00;
            16'd5369: data <= 8'hF8;
            16'd5370: data <= 8'h00;
            16'd5371: data <= 8'hF8;
            16'd5372: data <= 8'h00;
            16'd5373: data <= 8'hF8;
            16'd5374: data <= 8'h00;
            16'd5375: data <= 8'hF8;
            16'd5376: data <= 8'h00;
            16'd5377: data <= 8'hF8;
            16'd5378: data <= 8'h00;
            16'd5379: data <= 8'hF8;
            16'd5380: data <= 8'h00;
            16'd5381: data <= 8'hF8;
            16'd5382: data <= 8'h00;
            16'd5383: data <= 8'hF8;
            16'd5384: data <= 8'h00;
            16'd5385: data <= 8'hF8;
            16'd5386: data <= 8'h00;
            16'd5387: data <= 8'hF8;
            16'd5388: data <= 8'h00;
            16'd5389: data <= 8'hF8;
            16'd5390: data <= 8'h00;
            16'd5391: data <= 8'hF8;
            16'd5392: data <= 8'h00;
            16'd5393: data <= 8'hF8;
            16'd5394: data <= 8'h00;
            16'd5395: data <= 8'hF8;
            16'd5396: data <= 8'h00;
            16'd5397: data <= 8'hF8;
            16'd5398: data <= 8'h00;
            16'd5399: data <= 8'hF8;
            16'd5400: data <= 8'hFF;
            16'd5401: data <= 8'hFF;
            16'd5402: data <= 8'h00;
            16'd5403: data <= 8'hF8;
            16'd5404: data <= 8'h00;
            16'd5405: data <= 8'hF8;
            16'd5406: data <= 8'h00;
            16'd5407: data <= 8'hF8;
            16'd5408: data <= 8'h00;
            16'd5409: data <= 8'hF8;
            16'd5410: data <= 8'h00;
            16'd5411: data <= 8'hF8;
            16'd5412: data <= 8'h00;
            16'd5413: data <= 8'hF8;
            16'd5414: data <= 8'h00;
            16'd5415: data <= 8'hF8;
            16'd5416: data <= 8'h00;
            16'd5417: data <= 8'hF8;
            16'd5418: data <= 8'h00;
            16'd5419: data <= 8'hF8;
            16'd5420: data <= 8'h00;
            16'd5421: data <= 8'hF8;
            16'd5422: data <= 8'h00;
            16'd5423: data <= 8'hF8;
            16'd5424: data <= 8'h00;
            16'd5425: data <= 8'hF8;
            16'd5426: data <= 8'h00;
            16'd5427: data <= 8'hF8;
            16'd5428: data <= 8'h00;
            16'd5429: data <= 8'hF8;
            16'd5430: data <= 8'h00;
            16'd5431: data <= 8'hF8;
            16'd5432: data <= 8'h00;
            16'd5433: data <= 8'hF8;
            16'd5434: data <= 8'h00;
            16'd5435: data <= 8'hF8;
            16'd5436: data <= 8'h00;
            16'd5437: data <= 8'hF8;
            16'd5438: data <= 8'h00;
            16'd5439: data <= 8'hF8;
            16'd5440: data <= 8'hFF;
            16'd5441: data <= 8'hFF;
            16'd5442: data <= 8'h00;
            16'd5443: data <= 8'hF8;
            16'd5444: data <= 8'h00;
            16'd5445: data <= 8'hF8;
            16'd5446: data <= 8'h00;
            16'd5447: data <= 8'hF8;
            16'd5448: data <= 8'h00;
            16'd5449: data <= 8'hF8;
            16'd5450: data <= 8'h00;
            16'd5451: data <= 8'hF8;
            16'd5452: data <= 8'h00;
            16'd5453: data <= 8'hF8;
            16'd5454: data <= 8'h00;
            16'd5455: data <= 8'hF8;
            16'd5456: data <= 8'h00;
            16'd5457: data <= 8'hF8;
            16'd5458: data <= 8'h00;
            16'd5459: data <= 8'hF8;
            16'd5460: data <= 8'h00;
            16'd5461: data <= 8'hF8;
            16'd5462: data <= 8'h00;
            16'd5463: data <= 8'hF8;
            16'd5464: data <= 8'h00;
            16'd5465: data <= 8'hF8;
            16'd5466: data <= 8'h00;
            16'd5467: data <= 8'hF8;
            16'd5468: data <= 8'h00;
            16'd5469: data <= 8'hF8;
            16'd5470: data <= 8'h00;
            16'd5471: data <= 8'hF8;
            16'd5472: data <= 8'h00;
            16'd5473: data <= 8'hF8;
            16'd5474: data <= 8'h00;
            16'd5475: data <= 8'hF8;
            16'd5476: data <= 8'h00;
            16'd5477: data <= 8'hF8;
            16'd5478: data <= 8'h00;
            16'd5479: data <= 8'hF8;
            16'd5480: data <= 8'hFF;
            16'd5481: data <= 8'hFF;
            16'd5482: data <= 8'h00;
            16'd5483: data <= 8'hF8;
            16'd5484: data <= 8'h00;
            16'd5485: data <= 8'hF8;
            16'd5486: data <= 8'h00;
            16'd5487: data <= 8'hF8;
            16'd5488: data <= 8'h00;
            16'd5489: data <= 8'hF8;
            16'd5490: data <= 8'h00;
            16'd5491: data <= 8'hF8;
            16'd5492: data <= 8'h00;
            16'd5493: data <= 8'hF8;
            16'd5494: data <= 8'h00;
            16'd5495: data <= 8'hF8;
            16'd5496: data <= 8'h00;
            16'd5497: data <= 8'hF8;
            16'd5498: data <= 8'h00;
            16'd5499: data <= 8'hF8;
            16'd5500: data <= 8'h00;
            16'd5501: data <= 8'hF8;
            16'd5502: data <= 8'h00;
            16'd5503: data <= 8'hF8;
            16'd5504: data <= 8'h00;
            16'd5505: data <= 8'hF8;
            16'd5506: data <= 8'h00;
            16'd5507: data <= 8'hF8;
            16'd5508: data <= 8'h00;
            16'd5509: data <= 8'hF8;
            16'd5510: data <= 8'h00;
            16'd5511: data <= 8'hF8;
            16'd5512: data <= 8'h00;
            16'd5513: data <= 8'hF8;
            16'd5514: data <= 8'h00;
            16'd5515: data <= 8'hF8;
            16'd5516: data <= 8'h00;
            16'd5517: data <= 8'hF8;
            16'd5518: data <= 8'h00;
            16'd5519: data <= 8'hF8;
            16'd5520: data <= 8'hFF;
            16'd5521: data <= 8'hFF;
            16'd5522: data <= 8'h00;
            16'd5523: data <= 8'hF8;
            16'd5524: data <= 8'h00;
            16'd5525: data <= 8'hF8;
            16'd5526: data <= 8'h00;
            16'd5527: data <= 8'hF8;
            16'd5528: data <= 8'h00;
            16'd5529: data <= 8'hF8;
            16'd5530: data <= 8'h00;
            16'd5531: data <= 8'hF8;
            16'd5532: data <= 8'h00;
            16'd5533: data <= 8'hF8;
            16'd5534: data <= 8'h00;
            16'd5535: data <= 8'hF8;
            16'd5536: data <= 8'h00;
            16'd5537: data <= 8'hF8;
            16'd5538: data <= 8'h00;
            16'd5539: data <= 8'hF8;
            16'd5540: data <= 8'h00;
            16'd5541: data <= 8'hF8;
            16'd5542: data <= 8'h00;
            16'd5543: data <= 8'hF8;
            16'd5544: data <= 8'h00;
            16'd5545: data <= 8'hF8;
            16'd5546: data <= 8'h00;
            16'd5547: data <= 8'hF8;
            16'd5548: data <= 8'h00;
            16'd5549: data <= 8'hF8;
            16'd5550: data <= 8'h00;
            16'd5551: data <= 8'hF8;
            16'd5552: data <= 8'h00;
            16'd5553: data <= 8'hF8;
            16'd5554: data <= 8'h00;
            16'd5555: data <= 8'hF8;
            16'd5556: data <= 8'h00;
            16'd5557: data <= 8'hF8;
            16'd5558: data <= 8'h00;
            16'd5559: data <= 8'hF8;
            16'd5560: data <= 8'hFF;
            16'd5561: data <= 8'hFF;
            16'd5562: data <= 8'h00;
            16'd5563: data <= 8'hF8;
            16'd5564: data <= 8'h00;
            16'd5565: data <= 8'hF8;
            16'd5566: data <= 8'h00;
            16'd5567: data <= 8'hF8;
            16'd5568: data <= 8'h00;
            16'd5569: data <= 8'hF8;
            16'd5570: data <= 8'h00;
            16'd5571: data <= 8'hF8;
            16'd5572: data <= 8'h00;
            16'd5573: data <= 8'hF8;
            16'd5574: data <= 8'h00;
            16'd5575: data <= 8'hF8;
            16'd5576: data <= 8'h00;
            16'd5577: data <= 8'hF8;
            16'd5578: data <= 8'h00;
            16'd5579: data <= 8'hF8;
            16'd5580: data <= 8'h00;
            16'd5581: data <= 8'hF8;
            16'd5582: data <= 8'h00;
            16'd5583: data <= 8'hF8;
            16'd5584: data <= 8'h00;
            16'd5585: data <= 8'hF8;
            16'd5586: data <= 8'h00;
            16'd5587: data <= 8'hF8;
            16'd5588: data <= 8'h00;
            16'd5589: data <= 8'hF8;
            16'd5590: data <= 8'h00;
            16'd5591: data <= 8'hF8;
            16'd5592: data <= 8'h00;
            16'd5593: data <= 8'hF8;
            16'd5594: data <= 8'h00;
            16'd5595: data <= 8'hF8;
            16'd5596: data <= 8'h00;
            16'd5597: data <= 8'hF8;
            16'd5598: data <= 8'h00;
            16'd5599: data <= 8'hF8;
            16'd5600: data <= 8'hFF;
            16'd5601: data <= 8'hFF;
            16'd5602: data <= 8'h00;
            16'd5603: data <= 8'hF8;
            16'd5604: data <= 8'h00;
            16'd5605: data <= 8'hF8;
            16'd5606: data <= 8'h00;
            16'd5607: data <= 8'hF8;
            16'd5608: data <= 8'h00;
            16'd5609: data <= 8'hF8;
            16'd5610: data <= 8'h00;
            16'd5611: data <= 8'hF8;
            16'd5612: data <= 8'h00;
            16'd5613: data <= 8'hF8;
            16'd5614: data <= 8'h00;
            16'd5615: data <= 8'hF8;
            16'd5616: data <= 8'h00;
            16'd5617: data <= 8'hF8;
            16'd5618: data <= 8'h00;
            16'd5619: data <= 8'hF8;
            16'd5620: data <= 8'h00;
            16'd5621: data <= 8'hF8;
            16'd5622: data <= 8'h00;
            16'd5623: data <= 8'hF8;
            16'd5624: data <= 8'h00;
            16'd5625: data <= 8'hF8;
            16'd5626: data <= 8'h00;
            16'd5627: data <= 8'hF8;
            16'd5628: data <= 8'h00;
            16'd5629: data <= 8'hF8;
            16'd5630: data <= 8'h00;
            16'd5631: data <= 8'hF8;
            16'd5632: data <= 8'h00;
            16'd5633: data <= 8'hF8;
            16'd5634: data <= 8'h00;
            16'd5635: data <= 8'hF8;
            16'd5636: data <= 8'h00;
            16'd5637: data <= 8'hF8;
            16'd5638: data <= 8'h00;
            16'd5639: data <= 8'hF8;
            16'd5640: data <= 8'hFF;
            16'd5641: data <= 8'hFF;
            16'd5642: data <= 8'h00;
            16'd5643: data <= 8'hF8;
            16'd5644: data <= 8'h00;
            16'd5645: data <= 8'hF8;
            16'd5646: data <= 8'h00;
            16'd5647: data <= 8'hF8;
            16'd5648: data <= 8'h00;
            16'd5649: data <= 8'hF8;
            16'd5650: data <= 8'h00;
            16'd5651: data <= 8'hF8;
            16'd5652: data <= 8'h00;
            16'd5653: data <= 8'hF8;
            16'd5654: data <= 8'h00;
            16'd5655: data <= 8'hF8;
            16'd5656: data <= 8'h00;
            16'd5657: data <= 8'hF8;
            16'd5658: data <= 8'h00;
            16'd5659: data <= 8'hF8;
            16'd5660: data <= 8'h00;
            16'd5661: data <= 8'hF8;
            16'd5662: data <= 8'h00;
            16'd5663: data <= 8'hF8;
            16'd5664: data <= 8'h00;
            16'd5665: data <= 8'hF8;
            16'd5666: data <= 8'h00;
            16'd5667: data <= 8'hF8;
            16'd5668: data <= 8'h00;
            16'd5669: data <= 8'hF8;
            16'd5670: data <= 8'h00;
            16'd5671: data <= 8'hF8;
            16'd5672: data <= 8'h00;
            16'd5673: data <= 8'hF8;
            16'd5674: data <= 8'h00;
            16'd5675: data <= 8'hF8;
            16'd5676: data <= 8'h00;
            16'd5677: data <= 8'hF8;
            16'd5678: data <= 8'h00;
            16'd5679: data <= 8'hF8;
            16'd5680: data <= 8'hFF;
            16'd5681: data <= 8'hFF;
            16'd5682: data <= 8'h00;
            16'd5683: data <= 8'hF8;
            16'd5684: data <= 8'h00;
            16'd5685: data <= 8'hF8;
            16'd5686: data <= 8'h00;
            16'd5687: data <= 8'hF8;
            16'd5688: data <= 8'h00;
            16'd5689: data <= 8'hF8;
            16'd5690: data <= 8'h00;
            16'd5691: data <= 8'hF8;
            16'd5692: data <= 8'h00;
            16'd5693: data <= 8'hF8;
            16'd5694: data <= 8'h00;
            16'd5695: data <= 8'hF8;
            16'd5696: data <= 8'h00;
            16'd5697: data <= 8'hF8;
            16'd5698: data <= 8'h00;
            16'd5699: data <= 8'hF8;
            16'd5700: data <= 8'h00;
            16'd5701: data <= 8'hF8;
            16'd5702: data <= 8'h00;
            16'd5703: data <= 8'hF8;
            16'd5704: data <= 8'h00;
            16'd5705: data <= 8'hF8;
            16'd5706: data <= 8'h00;
            16'd5707: data <= 8'hF8;
            16'd5708: data <= 8'h00;
            16'd5709: data <= 8'hF8;
            16'd5710: data <= 8'h00;
            16'd5711: data <= 8'hF8;
            16'd5712: data <= 8'h00;
            16'd5713: data <= 8'hF8;
            16'd5714: data <= 8'h00;
            16'd5715: data <= 8'hF8;
            16'd5716: data <= 8'h00;
            16'd5717: data <= 8'hF8;
            16'd5718: data <= 8'h00;
            16'd5719: data <= 8'hF8;
            16'd5720: data <= 8'hFF;
            16'd5721: data <= 8'hFF;
            16'd5722: data <= 8'h00;
            16'd5723: data <= 8'hF8;
            16'd5724: data <= 8'h00;
            16'd5725: data <= 8'hF8;
            16'd5726: data <= 8'h00;
            16'd5727: data <= 8'hF8;
            16'd5728: data <= 8'h00;
            16'd5729: data <= 8'hF8;
            16'd5730: data <= 8'h00;
            16'd5731: data <= 8'hF8;
            16'd5732: data <= 8'h00;
            16'd5733: data <= 8'hF8;
            16'd5734: data <= 8'h00;
            16'd5735: data <= 8'hF8;
            16'd5736: data <= 8'h00;
            16'd5737: data <= 8'hF8;
            16'd5738: data <= 8'h00;
            16'd5739: data <= 8'hF8;
            16'd5740: data <= 8'h00;
            16'd5741: data <= 8'hF8;
            16'd5742: data <= 8'h00;
            16'd5743: data <= 8'hF8;
            16'd5744: data <= 8'h00;
            16'd5745: data <= 8'hF8;
            16'd5746: data <= 8'h00;
            16'd5747: data <= 8'hF8;
            16'd5748: data <= 8'h00;
            16'd5749: data <= 8'hF8;
            16'd5750: data <= 8'h00;
            16'd5751: data <= 8'hF8;
            16'd5752: data <= 8'h00;
            16'd5753: data <= 8'hF8;
            16'd5754: data <= 8'h00;
            16'd5755: data <= 8'hF8;
            16'd5756: data <= 8'h00;
            16'd5757: data <= 8'hF8;
            16'd5758: data <= 8'h00;
            16'd5759: data <= 8'hF8;
            16'd5760: data <= 8'hFF;
            16'd5761: data <= 8'hFF;
            16'd5762: data <= 8'h00;
            16'd5763: data <= 8'hF8;
            16'd5764: data <= 8'h00;
            16'd5765: data <= 8'hF8;
            16'd5766: data <= 8'h00;
            16'd5767: data <= 8'hF8;
            16'd5768: data <= 8'h00;
            16'd5769: data <= 8'hF8;
            16'd5770: data <= 8'h00;
            16'd5771: data <= 8'hF8;
            16'd5772: data <= 8'h00;
            16'd5773: data <= 8'hF8;
            16'd5774: data <= 8'h00;
            16'd5775: data <= 8'hF8;
            16'd5776: data <= 8'h00;
            16'd5777: data <= 8'hF8;
            16'd5778: data <= 8'h00;
            16'd5779: data <= 8'hF8;
            16'd5780: data <= 8'h00;
            16'd5781: data <= 8'hF8;
            16'd5782: data <= 8'h00;
            16'd5783: data <= 8'hF8;
            16'd5784: data <= 8'h00;
            16'd5785: data <= 8'hF8;
            16'd5786: data <= 8'h00;
            16'd5787: data <= 8'hF8;
            16'd5788: data <= 8'h00;
            16'd5789: data <= 8'hF8;
            16'd5790: data <= 8'h00;
            16'd5791: data <= 8'hF8;
            16'd5792: data <= 8'h00;
            16'd5793: data <= 8'hF8;
            16'd5794: data <= 8'h00;
            16'd5795: data <= 8'hF8;
            16'd5796: data <= 8'h00;
            16'd5797: data <= 8'hF8;
            16'd5798: data <= 8'h00;
            16'd5799: data <= 8'hF8;
            16'd5800: data <= 8'hFF;
            16'd5801: data <= 8'hFF;
            16'd5802: data <= 8'h00;
            16'd5803: data <= 8'hF8;
            16'd5804: data <= 8'h00;
            16'd5805: data <= 8'hF8;
            16'd5806: data <= 8'h00;
            16'd5807: data <= 8'hF8;
            16'd5808: data <= 8'h00;
            16'd5809: data <= 8'hF8;
            16'd5810: data <= 8'h00;
            16'd5811: data <= 8'hF8;
            16'd5812: data <= 8'h00;
            16'd5813: data <= 8'hF8;
            16'd5814: data <= 8'h00;
            16'd5815: data <= 8'hF8;
            16'd5816: data <= 8'h00;
            16'd5817: data <= 8'hF8;
            16'd5818: data <= 8'h00;
            16'd5819: data <= 8'hF8;
            16'd5820: data <= 8'h00;
            16'd5821: data <= 8'hF8;
            16'd5822: data <= 8'h00;
            16'd5823: data <= 8'hF8;
            16'd5824: data <= 8'h00;
            16'd5825: data <= 8'hF8;
            16'd5826: data <= 8'h00;
            16'd5827: data <= 8'hF8;
            16'd5828: data <= 8'h00;
            16'd5829: data <= 8'hF8;
            16'd5830: data <= 8'h00;
            16'd5831: data <= 8'hF8;
            16'd5832: data <= 8'h00;
            16'd5833: data <= 8'hF8;
            16'd5834: data <= 8'h00;
            16'd5835: data <= 8'hF8;
            16'd5836: data <= 8'h00;
            16'd5837: data <= 8'hF8;
            16'd5838: data <= 8'h00;
            16'd5839: data <= 8'hF8;
            16'd5840: data <= 8'hFF;
            16'd5841: data <= 8'hFF;
            16'd5842: data <= 8'h00;
            16'd5843: data <= 8'hF8;
            16'd5844: data <= 8'h00;
            16'd5845: data <= 8'hF8;
            16'd5846: data <= 8'h00;
            16'd5847: data <= 8'hF8;
            16'd5848: data <= 8'h00;
            16'd5849: data <= 8'hF8;
            16'd5850: data <= 8'h00;
            16'd5851: data <= 8'hF8;
            16'd5852: data <= 8'h00;
            16'd5853: data <= 8'hF8;
            16'd5854: data <= 8'h00;
            16'd5855: data <= 8'hF8;
            16'd5856: data <= 8'h00;
            16'd5857: data <= 8'hF8;
            16'd5858: data <= 8'h00;
            16'd5859: data <= 8'hF8;
            16'd5860: data <= 8'h00;
            16'd5861: data <= 8'hF8;
            16'd5862: data <= 8'h00;
            16'd5863: data <= 8'hF8;
            16'd5864: data <= 8'h00;
            16'd5865: data <= 8'hF8;
            16'd5866: data <= 8'h00;
            16'd5867: data <= 8'hF8;
            16'd5868: data <= 8'h00;
            16'd5869: data <= 8'hF8;
            16'd5870: data <= 8'h00;
            16'd5871: data <= 8'hF8;
            16'd5872: data <= 8'h00;
            16'd5873: data <= 8'hF8;
            16'd5874: data <= 8'h00;
            16'd5875: data <= 8'hF8;
            16'd5876: data <= 8'h00;
            16'd5877: data <= 8'hF8;
            16'd5878: data <= 8'h00;
            16'd5879: data <= 8'hF8;
            16'd5880: data <= 8'hFF;
            16'd5881: data <= 8'hFF;
            16'd5882: data <= 8'h00;
            16'd5883: data <= 8'hF8;
            16'd5884: data <= 8'h00;
            16'd5885: data <= 8'hF8;
            16'd5886: data <= 8'h00;
            16'd5887: data <= 8'hF8;
            16'd5888: data <= 8'h00;
            16'd5889: data <= 8'hF8;
            16'd5890: data <= 8'h00;
            16'd5891: data <= 8'hF8;
            16'd5892: data <= 8'h00;
            16'd5893: data <= 8'hF8;
            16'd5894: data <= 8'h00;
            16'd5895: data <= 8'hF8;
            16'd5896: data <= 8'h00;
            16'd5897: data <= 8'hF8;
            16'd5898: data <= 8'h00;
            16'd5899: data <= 8'hF8;
            16'd5900: data <= 8'h00;
            16'd5901: data <= 8'hF8;
            16'd5902: data <= 8'h00;
            16'd5903: data <= 8'hF8;
            16'd5904: data <= 8'h00;
            16'd5905: data <= 8'hF8;
            16'd5906: data <= 8'h00;
            16'd5907: data <= 8'hF8;
            16'd5908: data <= 8'h00;
            16'd5909: data <= 8'hF8;
            16'd5910: data <= 8'h00;
            16'd5911: data <= 8'hF8;
            16'd5912: data <= 8'h00;
            16'd5913: data <= 8'hF8;
            16'd5914: data <= 8'h00;
            16'd5915: data <= 8'hF8;
            16'd5916: data <= 8'h00;
            16'd5917: data <= 8'hF8;
            16'd5918: data <= 8'h00;
            16'd5919: data <= 8'hF8;
            16'd5920: data <= 8'hFF;
            16'd5921: data <= 8'hFF;
            16'd5922: data <= 8'h00;
            16'd5923: data <= 8'hF8;
            16'd5924: data <= 8'h00;
            16'd5925: data <= 8'hF8;
            16'd5926: data <= 8'h00;
            16'd5927: data <= 8'hF8;
            16'd5928: data <= 8'h00;
            16'd5929: data <= 8'hF8;
            16'd5930: data <= 8'h00;
            16'd5931: data <= 8'hF8;
            16'd5932: data <= 8'h00;
            16'd5933: data <= 8'hF8;
            16'd5934: data <= 8'h00;
            16'd5935: data <= 8'hF8;
            16'd5936: data <= 8'h00;
            16'd5937: data <= 8'hF8;
            16'd5938: data <= 8'h00;
            16'd5939: data <= 8'hF8;
            16'd5940: data <= 8'h00;
            16'd5941: data <= 8'hF8;
            16'd5942: data <= 8'h00;
            16'd5943: data <= 8'hF8;
            16'd5944: data <= 8'h00;
            16'd5945: data <= 8'hF8;
            16'd5946: data <= 8'h00;
            16'd5947: data <= 8'hF8;
            16'd5948: data <= 8'h00;
            16'd5949: data <= 8'hF8;
            16'd5950: data <= 8'h00;
            16'd5951: data <= 8'hF8;
            16'd5952: data <= 8'h00;
            16'd5953: data <= 8'hF8;
            16'd5954: data <= 8'h00;
            16'd5955: data <= 8'hF8;
            16'd5956: data <= 8'h00;
            16'd5957: data <= 8'hF8;
            16'd5958: data <= 8'h00;
            16'd5959: data <= 8'hF8;
            16'd5960: data <= 8'hFF;
            16'd5961: data <= 8'hFF;
            16'd5962: data <= 8'h00;
            16'd5963: data <= 8'hF8;
            16'd5964: data <= 8'h00;
            16'd5965: data <= 8'hF8;
            16'd5966: data <= 8'h00;
            16'd5967: data <= 8'hF8;
            16'd5968: data <= 8'h00;
            16'd5969: data <= 8'hF8;
            16'd5970: data <= 8'h00;
            16'd5971: data <= 8'hF8;
            16'd5972: data <= 8'h00;
            16'd5973: data <= 8'hF8;
            16'd5974: data <= 8'h00;
            16'd5975: data <= 8'hF8;
            16'd5976: data <= 8'h00;
            16'd5977: data <= 8'hF8;
            16'd5978: data <= 8'h00;
            16'd5979: data <= 8'hF8;
            16'd5980: data <= 8'h00;
            16'd5981: data <= 8'hF8;
            16'd5982: data <= 8'h00;
            16'd5983: data <= 8'hF8;
            16'd5984: data <= 8'h00;
            16'd5985: data <= 8'hF8;
            16'd5986: data <= 8'h00;
            16'd5987: data <= 8'hF8;
            16'd5988: data <= 8'h00;
            16'd5989: data <= 8'hF8;
            16'd5990: data <= 8'h00;
            16'd5991: data <= 8'hF8;
            16'd5992: data <= 8'h00;
            16'd5993: data <= 8'hF8;
            16'd5994: data <= 8'h00;
            16'd5995: data <= 8'hF8;
            16'd5996: data <= 8'h00;
            16'd5997: data <= 8'hF8;
            16'd5998: data <= 8'h00;
            16'd5999: data <= 8'hF8;
            16'd6000: data <= 8'hFF;
            16'd6001: data <= 8'hFF;
            16'd6002: data <= 8'h00;
            16'd6003: data <= 8'hF8;
            16'd6004: data <= 8'h00;
            16'd6005: data <= 8'hF8;
            16'd6006: data <= 8'h00;
            16'd6007: data <= 8'hF8;
            16'd6008: data <= 8'h00;
            16'd6009: data <= 8'hF8;
            16'd6010: data <= 8'h00;
            16'd6011: data <= 8'hF8;
            16'd6012: data <= 8'h00;
            16'd6013: data <= 8'hF8;
            16'd6014: data <= 8'h00;
            16'd6015: data <= 8'hF8;
            16'd6016: data <= 8'h00;
            16'd6017: data <= 8'hF8;
            16'd6018: data <= 8'h00;
            16'd6019: data <= 8'hF8;
            16'd6020: data <= 8'h00;
            16'd6021: data <= 8'hF8;
            16'd6022: data <= 8'h00;
            16'd6023: data <= 8'hF8;
            16'd6024: data <= 8'h00;
            16'd6025: data <= 8'hF8;
            16'd6026: data <= 8'h00;
            16'd6027: data <= 8'hF8;
            16'd6028: data <= 8'h00;
            16'd6029: data <= 8'hF8;
            16'd6030: data <= 8'h00;
            16'd6031: data <= 8'hF8;
            16'd6032: data <= 8'h00;
            16'd6033: data <= 8'hF8;
            16'd6034: data <= 8'h00;
            16'd6035: data <= 8'hF8;
            16'd6036: data <= 8'h00;
            16'd6037: data <= 8'hF8;
            16'd6038: data <= 8'h00;
            16'd6039: data <= 8'hF8;
            16'd6040: data <= 8'hFF;
            16'd6041: data <= 8'hFF;
            16'd6042: data <= 8'h00;
            16'd6043: data <= 8'hF8;
            16'd6044: data <= 8'h00;
            16'd6045: data <= 8'hF8;
            16'd6046: data <= 8'h00;
            16'd6047: data <= 8'hF8;
            16'd6048: data <= 8'h00;
            16'd6049: data <= 8'hF8;
            16'd6050: data <= 8'h00;
            16'd6051: data <= 8'hF8;
            16'd6052: data <= 8'h00;
            16'd6053: data <= 8'hF8;
            16'd6054: data <= 8'h00;
            16'd6055: data <= 8'hF8;
            16'd6056: data <= 8'h00;
            16'd6057: data <= 8'hF8;
            16'd6058: data <= 8'h00;
            16'd6059: data <= 8'hF8;
            16'd6060: data <= 8'h00;
            16'd6061: data <= 8'hF8;
            16'd6062: data <= 8'h00;
            16'd6063: data <= 8'hF8;
            16'd6064: data <= 8'h00;
            16'd6065: data <= 8'hF8;
            16'd6066: data <= 8'h00;
            16'd6067: data <= 8'hF8;
            16'd6068: data <= 8'h00;
            16'd6069: data <= 8'hF8;
            16'd6070: data <= 8'h00;
            16'd6071: data <= 8'hF8;
            16'd6072: data <= 8'h00;
            16'd6073: data <= 8'hF8;
            16'd6074: data <= 8'h00;
            16'd6075: data <= 8'hF8;
            16'd6076: data <= 8'h00;
            16'd6077: data <= 8'hF8;
            16'd6078: data <= 8'h00;
            16'd6079: data <= 8'hF8;
            16'd6080: data <= 8'hFF;
            16'd6081: data <= 8'hFF;
            16'd6082: data <= 8'h00;
            16'd6083: data <= 8'hF8;
            16'd6084: data <= 8'h00;
            16'd6085: data <= 8'hF8;
            16'd6086: data <= 8'h00;
            16'd6087: data <= 8'hF8;
            16'd6088: data <= 8'h00;
            16'd6089: data <= 8'hF8;
            16'd6090: data <= 8'h00;
            16'd6091: data <= 8'hF8;
            16'd6092: data <= 8'h00;
            16'd6093: data <= 8'hF8;
            16'd6094: data <= 8'h00;
            16'd6095: data <= 8'hF8;
            16'd6096: data <= 8'h00;
            16'd6097: data <= 8'hF8;
            16'd6098: data <= 8'h00;
            16'd6099: data <= 8'hF8;
            16'd6100: data <= 8'h00;
            16'd6101: data <= 8'hF8;
            16'd6102: data <= 8'h00;
            16'd6103: data <= 8'hF8;
            16'd6104: data <= 8'h00;
            16'd6105: data <= 8'hF8;
            16'd6106: data <= 8'h00;
            16'd6107: data <= 8'hF8;
            16'd6108: data <= 8'h00;
            16'd6109: data <= 8'hF8;
            16'd6110: data <= 8'h00;
            16'd6111: data <= 8'hF8;
            16'd6112: data <= 8'h00;
            16'd6113: data <= 8'hF8;
            16'd6114: data <= 8'h00;
            16'd6115: data <= 8'hF8;
            16'd6116: data <= 8'h00;
            16'd6117: data <= 8'hF8;
            16'd6118: data <= 8'h00;
            16'd6119: data <= 8'hF8;
            16'd6120: data <= 8'hFF;
            16'd6121: data <= 8'hFF;
            16'd6122: data <= 8'h00;
            16'd6123: data <= 8'hF8;
            16'd6124: data <= 8'h00;
            16'd6125: data <= 8'hF8;
            16'd6126: data <= 8'h00;
            16'd6127: data <= 8'hF8;
            16'd6128: data <= 8'h00;
            16'd6129: data <= 8'hF8;
            16'd6130: data <= 8'h00;
            16'd6131: data <= 8'hF8;
            16'd6132: data <= 8'h00;
            16'd6133: data <= 8'hF8;
            16'd6134: data <= 8'h00;
            16'd6135: data <= 8'hF8;
            16'd6136: data <= 8'h00;
            16'd6137: data <= 8'hF8;
            16'd6138: data <= 8'h00;
            16'd6139: data <= 8'hF8;
            16'd6140: data <= 8'h00;
            16'd6141: data <= 8'hF8;
            16'd6142: data <= 8'h00;
            16'd6143: data <= 8'hF8;
            16'd6144: data <= 8'h00;
            16'd6145: data <= 8'hF8;
            16'd6146: data <= 8'h00;
            16'd6147: data <= 8'hF8;
            16'd6148: data <= 8'h00;
            16'd6149: data <= 8'hF8;
            16'd6150: data <= 8'h00;
            16'd6151: data <= 8'hF8;
            16'd6152: data <= 8'h00;
            16'd6153: data <= 8'hF8;
            16'd6154: data <= 8'h00;
            16'd6155: data <= 8'hF8;
            16'd6156: data <= 8'h00;
            16'd6157: data <= 8'hF8;
            16'd6158: data <= 8'h00;
            16'd6159: data <= 8'hF8;
            16'd6160: data <= 8'hFF;
            16'd6161: data <= 8'hFF;
            16'd6162: data <= 8'h00;
            16'd6163: data <= 8'hF8;
            16'd6164: data <= 8'h00;
            16'd6165: data <= 8'hF8;
            16'd6166: data <= 8'h00;
            16'd6167: data <= 8'hF8;
            16'd6168: data <= 8'h00;
            16'd6169: data <= 8'hF8;
            16'd6170: data <= 8'h00;
            16'd6171: data <= 8'hF8;
            16'd6172: data <= 8'h00;
            16'd6173: data <= 8'hF8;
            16'd6174: data <= 8'h00;
            16'd6175: data <= 8'hF8;
            16'd6176: data <= 8'h00;
            16'd6177: data <= 8'hF8;
            16'd6178: data <= 8'h00;
            16'd6179: data <= 8'hF8;
            16'd6180: data <= 8'h00;
            16'd6181: data <= 8'hF8;
            16'd6182: data <= 8'h00;
            16'd6183: data <= 8'hF8;
            16'd6184: data <= 8'h00;
            16'd6185: data <= 8'hF8;
            16'd6186: data <= 8'h00;
            16'd6187: data <= 8'hF8;
            16'd6188: data <= 8'h00;
            16'd6189: data <= 8'hF8;
            16'd6190: data <= 8'h00;
            16'd6191: data <= 8'hF8;
            16'd6192: data <= 8'h00;
            16'd6193: data <= 8'hF8;
            16'd6194: data <= 8'h00;
            16'd6195: data <= 8'hF8;
            16'd6196: data <= 8'h00;
            16'd6197: data <= 8'hF8;
            16'd6198: data <= 8'h00;
            16'd6199: data <= 8'hF8;
            16'd6200: data <= 8'hFF;
            16'd6201: data <= 8'hFF;
            16'd6202: data <= 8'h00;
            16'd6203: data <= 8'hF8;
            16'd6204: data <= 8'h00;
            16'd6205: data <= 8'hF8;
            16'd6206: data <= 8'h00;
            16'd6207: data <= 8'hF8;
            16'd6208: data <= 8'h00;
            16'd6209: data <= 8'hF8;
            16'd6210: data <= 8'h00;
            16'd6211: data <= 8'hF8;
            16'd6212: data <= 8'h00;
            16'd6213: data <= 8'hF8;
            16'd6214: data <= 8'h00;
            16'd6215: data <= 8'hF8;
            16'd6216: data <= 8'h00;
            16'd6217: data <= 8'hF8;
            16'd6218: data <= 8'h00;
            16'd6219: data <= 8'hF8;
            16'd6220: data <= 8'h00;
            16'd6221: data <= 8'hF8;
            16'd6222: data <= 8'h00;
            16'd6223: data <= 8'hF8;
            16'd6224: data <= 8'h00;
            16'd6225: data <= 8'hF8;
            16'd6226: data <= 8'h00;
            16'd6227: data <= 8'hF8;
            16'd6228: data <= 8'h00;
            16'd6229: data <= 8'hF8;
            16'd6230: data <= 8'h00;
            16'd6231: data <= 8'hF8;
            16'd6232: data <= 8'h00;
            16'd6233: data <= 8'hF8;
            16'd6234: data <= 8'h00;
            16'd6235: data <= 8'hF8;
            16'd6236: data <= 8'h00;
            16'd6237: data <= 8'hF8;
            16'd6238: data <= 8'h00;
            16'd6239: data <= 8'hF8;
            16'd6240: data <= 8'hFF;
            16'd6241: data <= 8'hFF;
            16'd6242: data <= 8'h00;
            16'd6243: data <= 8'hF8;
            16'd6244: data <= 8'h00;
            16'd6245: data <= 8'hF8;
            16'd6246: data <= 8'h00;
            16'd6247: data <= 8'hF8;
            16'd6248: data <= 8'h00;
            16'd6249: data <= 8'hF8;
            16'd6250: data <= 8'h00;
            16'd6251: data <= 8'hF8;
            16'd6252: data <= 8'h00;
            16'd6253: data <= 8'hF8;
            16'd6254: data <= 8'h00;
            16'd6255: data <= 8'hF8;
            16'd6256: data <= 8'h00;
            16'd6257: data <= 8'hF8;
            16'd6258: data <= 8'h00;
            16'd6259: data <= 8'hF8;
            16'd6260: data <= 8'h00;
            16'd6261: data <= 8'hF8;
            16'd6262: data <= 8'h00;
            16'd6263: data <= 8'hF8;
            16'd6264: data <= 8'h00;
            16'd6265: data <= 8'hF8;
            16'd6266: data <= 8'h00;
            16'd6267: data <= 8'hF8;
            16'd6268: data <= 8'h00;
            16'd6269: data <= 8'hF8;
            16'd6270: data <= 8'h00;
            16'd6271: data <= 8'hF8;
            16'd6272: data <= 8'h00;
            16'd6273: data <= 8'hF8;
            16'd6274: data <= 8'h00;
            16'd6275: data <= 8'hF8;
            16'd6276: data <= 8'h00;
            16'd6277: data <= 8'hF8;
            16'd6278: data <= 8'h00;
            16'd6279: data <= 8'hF8;
            16'd6280: data <= 8'hFF;
            16'd6281: data <= 8'hFF;
            16'd6282: data <= 8'h00;
            16'd6283: data <= 8'hF8;
            16'd6284: data <= 8'h00;
            16'd6285: data <= 8'hF8;
            16'd6286: data <= 8'h00;
            16'd6287: data <= 8'hF8;
            16'd6288: data <= 8'h00;
            16'd6289: data <= 8'hF8;
            16'd6290: data <= 8'h00;
            16'd6291: data <= 8'hF8;
            16'd6292: data <= 8'h00;
            16'd6293: data <= 8'hF8;
            16'd6294: data <= 8'h00;
            16'd6295: data <= 8'hF8;
            16'd6296: data <= 8'h00;
            16'd6297: data <= 8'hF8;
            16'd6298: data <= 8'h00;
            16'd6299: data <= 8'hF8;
            16'd6300: data <= 8'h00;
            16'd6301: data <= 8'hF8;
            16'd6302: data <= 8'h00;
            16'd6303: data <= 8'hF8;
            16'd6304: data <= 8'h00;
            16'd6305: data <= 8'hF8;
            16'd6306: data <= 8'h00;
            16'd6307: data <= 8'hF8;
            16'd6308: data <= 8'h00;
            16'd6309: data <= 8'hF8;
            16'd6310: data <= 8'h00;
            16'd6311: data <= 8'hF8;
            16'd6312: data <= 8'h00;
            16'd6313: data <= 8'hF8;
            16'd6314: data <= 8'h00;
            16'd6315: data <= 8'hF8;
            16'd6316: data <= 8'h00;
            16'd6317: data <= 8'hF8;
            16'd6318: data <= 8'h00;
            16'd6319: data <= 8'hF8;
            16'd6320: data <= 8'hFF;
            16'd6321: data <= 8'hFF;
            16'd6322: data <= 8'h00;
            16'd6323: data <= 8'hF8;
            16'd6324: data <= 8'h00;
            16'd6325: data <= 8'hF8;
            16'd6326: data <= 8'h00;
            16'd6327: data <= 8'hF8;
            16'd6328: data <= 8'h00;
            16'd6329: data <= 8'hF8;
            16'd6330: data <= 8'h00;
            16'd6331: data <= 8'hF8;
            16'd6332: data <= 8'h00;
            16'd6333: data <= 8'hF8;
            16'd6334: data <= 8'h00;
            16'd6335: data <= 8'hF8;
            16'd6336: data <= 8'h00;
            16'd6337: data <= 8'hF8;
            16'd6338: data <= 8'h00;
            16'd6339: data <= 8'hF8;
            16'd6340: data <= 8'h00;
            16'd6341: data <= 8'hF8;
            16'd6342: data <= 8'h00;
            16'd6343: data <= 8'hF8;
            16'd6344: data <= 8'h00;
            16'd6345: data <= 8'hF8;
            16'd6346: data <= 8'h00;
            16'd6347: data <= 8'hF8;
            16'd6348: data <= 8'h00;
            16'd6349: data <= 8'hF8;
            16'd6350: data <= 8'h00;
            16'd6351: data <= 8'hF8;
            16'd6352: data <= 8'h00;
            16'd6353: data <= 8'hF8;
            16'd6354: data <= 8'h00;
            16'd6355: data <= 8'hF8;
            16'd6356: data <= 8'h00;
            16'd6357: data <= 8'hF8;
            16'd6358: data <= 8'h00;
            16'd6359: data <= 8'hF8;
            16'd6360: data <= 8'hFF;
            16'd6361: data <= 8'hFF;
            16'd6362: data <= 8'h00;
            16'd6363: data <= 8'hF8;
            16'd6364: data <= 8'h00;
            16'd6365: data <= 8'hF8;
            16'd6366: data <= 8'h00;
            16'd6367: data <= 8'hF8;
            16'd6368: data <= 8'h00;
            16'd6369: data <= 8'hF8;
            16'd6370: data <= 8'h00;
            16'd6371: data <= 8'hF8;
            16'd6372: data <= 8'h00;
            16'd6373: data <= 8'hF8;
            16'd6374: data <= 8'h00;
            16'd6375: data <= 8'hF8;
            16'd6376: data <= 8'h00;
            16'd6377: data <= 8'hF8;
            16'd6378: data <= 8'h00;
            16'd6379: data <= 8'hF8;
            16'd6380: data <= 8'h00;
            16'd6381: data <= 8'hF8;
            16'd6382: data <= 8'h00;
            16'd6383: data <= 8'hF8;
            16'd6384: data <= 8'h00;
            16'd6385: data <= 8'hF8;
            16'd6386: data <= 8'h00;
            16'd6387: data <= 8'hF8;
            16'd6388: data <= 8'h00;
            16'd6389: data <= 8'hF8;
            16'd6390: data <= 8'h00;
            16'd6391: data <= 8'hF8;
            16'd6392: data <= 8'h00;
            16'd6393: data <= 8'hF8;
            16'd6394: data <= 8'h00;
            16'd6395: data <= 8'hF8;
            16'd6396: data <= 8'h00;
            16'd6397: data <= 8'hF8;
            16'd6398: data <= 8'h00;
            16'd6399: data <= 8'hF8;
            16'd6400: data <= 8'hFF;
            16'd6401: data <= 8'hFF;
            16'd6402: data <= 8'h00;
            16'd6403: data <= 8'hF8;
            16'd6404: data <= 8'h00;
            16'd6405: data <= 8'hF8;
            16'd6406: data <= 8'h00;
            16'd6407: data <= 8'hF8;
            16'd6408: data <= 8'h00;
            16'd6409: data <= 8'hF8;
            16'd6410: data <= 8'h00;
            16'd6411: data <= 8'hF8;
            16'd6412: data <= 8'h00;
            16'd6413: data <= 8'hF8;
            16'd6414: data <= 8'h00;
            16'd6415: data <= 8'hF8;
            16'd6416: data <= 8'h00;
            16'd6417: data <= 8'hF8;
            16'd6418: data <= 8'h00;
            16'd6419: data <= 8'hF8;
            16'd6420: data <= 8'h00;
            16'd6421: data <= 8'hF8;
            16'd6422: data <= 8'h00;
            16'd6423: data <= 8'hF8;
            16'd6424: data <= 8'h00;
            16'd6425: data <= 8'hF8;
            16'd6426: data <= 8'h00;
            16'd6427: data <= 8'hF8;
            16'd6428: data <= 8'h00;
            16'd6429: data <= 8'hF8;
            16'd6430: data <= 8'h00;
            16'd6431: data <= 8'hF8;
            16'd6432: data <= 8'h00;
            16'd6433: data <= 8'hF8;
            16'd6434: data <= 8'h00;
            16'd6435: data <= 8'hF8;
            16'd6436: data <= 8'h00;
            16'd6437: data <= 8'hF8;
            16'd6438: data <= 8'h00;
            16'd6439: data <= 8'hF8;
            16'd6440: data <= 8'hFF;
            16'd6441: data <= 8'hFF;
            16'd6442: data <= 8'h00;
            16'd6443: data <= 8'hF8;
            16'd6444: data <= 8'h00;
            16'd6445: data <= 8'hF8;
            16'd6446: data <= 8'h00;
            16'd6447: data <= 8'hF8;
            16'd6448: data <= 8'h00;
            16'd6449: data <= 8'hF8;
            16'd6450: data <= 8'h00;
            16'd6451: data <= 8'hF8;
            16'd6452: data <= 8'h00;
            16'd6453: data <= 8'hF8;
            16'd6454: data <= 8'h00;
            16'd6455: data <= 8'hF8;
            16'd6456: data <= 8'h00;
            16'd6457: data <= 8'hF8;
            16'd6458: data <= 8'h00;
            16'd6459: data <= 8'hF8;
            16'd6460: data <= 8'h00;
            16'd6461: data <= 8'hF8;
            16'd6462: data <= 8'h00;
            16'd6463: data <= 8'hF8;
            16'd6464: data <= 8'h00;
            16'd6465: data <= 8'hF8;
            16'd6466: data <= 8'h00;
            16'd6467: data <= 8'hF8;
            16'd6468: data <= 8'h00;
            16'd6469: data <= 8'hF8;
            16'd6470: data <= 8'h00;
            16'd6471: data <= 8'hF8;
            16'd6472: data <= 8'h00;
            16'd6473: data <= 8'hF8;
            16'd6474: data <= 8'h00;
            16'd6475: data <= 8'hF8;
            16'd6476: data <= 8'h00;
            16'd6477: data <= 8'hF8;
            16'd6478: data <= 8'h00;
            16'd6479: data <= 8'hF8;
            16'd6480: data <= 8'hFF;
            16'd6481: data <= 8'hFF;
            16'd6482: data <= 8'h00;
            16'd6483: data <= 8'hF8;
            16'd6484: data <= 8'h00;
            16'd6485: data <= 8'hF8;
            16'd6486: data <= 8'h00;
            16'd6487: data <= 8'hF8;
            16'd6488: data <= 8'h00;
            16'd6489: data <= 8'hF8;
            16'd6490: data <= 8'h00;
            16'd6491: data <= 8'hF8;
            16'd6492: data <= 8'h00;
            16'd6493: data <= 8'hF8;
            16'd6494: data <= 8'h00;
            16'd6495: data <= 8'hF8;
            16'd6496: data <= 8'h00;
            16'd6497: data <= 8'hF8;
            16'd6498: data <= 8'h00;
            16'd6499: data <= 8'hF8;
            16'd6500: data <= 8'h00;
            16'd6501: data <= 8'hF8;
            16'd6502: data <= 8'h00;
            16'd6503: data <= 8'hF8;
            16'd6504: data <= 8'h00;
            16'd6505: data <= 8'hF8;
            16'd6506: data <= 8'h00;
            16'd6507: data <= 8'hF8;
            16'd6508: data <= 8'h00;
            16'd6509: data <= 8'hF8;
            16'd6510: data <= 8'h00;
            16'd6511: data <= 8'hF8;
            16'd6512: data <= 8'h00;
            16'd6513: data <= 8'hF8;
            16'd6514: data <= 8'h00;
            16'd6515: data <= 8'hF8;
            16'd6516: data <= 8'h00;
            16'd6517: data <= 8'hF8;
            16'd6518: data <= 8'h00;
            16'd6519: data <= 8'hF8;
            16'd6520: data <= 8'hFF;
            16'd6521: data <= 8'hFF;
            16'd6522: data <= 8'h00;
            16'd6523: data <= 8'hF8;
            16'd6524: data <= 8'h00;
            16'd6525: data <= 8'hF8;
            16'd6526: data <= 8'h00;
            16'd6527: data <= 8'hF8;
            16'd6528: data <= 8'h00;
            16'd6529: data <= 8'hF8;
            16'd6530: data <= 8'h00;
            16'd6531: data <= 8'hF8;
            16'd6532: data <= 8'h00;
            16'd6533: data <= 8'hF8;
            16'd6534: data <= 8'h00;
            16'd6535: data <= 8'hF8;
            16'd6536: data <= 8'h00;
            16'd6537: data <= 8'hF8;
            16'd6538: data <= 8'h00;
            16'd6539: data <= 8'hF8;
            16'd6540: data <= 8'h00;
            16'd6541: data <= 8'hF8;
            16'd6542: data <= 8'h00;
            16'd6543: data <= 8'hF8;
            16'd6544: data <= 8'h00;
            16'd6545: data <= 8'hF8;
            16'd6546: data <= 8'h00;
            16'd6547: data <= 8'hF8;
            16'd6548: data <= 8'h00;
            16'd6549: data <= 8'hF8;
            16'd6550: data <= 8'h00;
            16'd6551: data <= 8'hF8;
            16'd6552: data <= 8'h00;
            16'd6553: data <= 8'hF8;
            16'd6554: data <= 8'h00;
            16'd6555: data <= 8'hF8;
            16'd6556: data <= 8'h00;
            16'd6557: data <= 8'hF8;
            16'd6558: data <= 8'h00;
            16'd6559: data <= 8'hF8;
            16'd6560: data <= 8'hFF;
            16'd6561: data <= 8'hFF;
            16'd6562: data <= 8'h00;
            16'd6563: data <= 8'hF8;
            16'd6564: data <= 8'h00;
            16'd6565: data <= 8'hF8;
            16'd6566: data <= 8'h00;
            16'd6567: data <= 8'hF8;
            16'd6568: data <= 8'h00;
            16'd6569: data <= 8'hF8;
            16'd6570: data <= 8'h00;
            16'd6571: data <= 8'hF8;
            16'd6572: data <= 8'h00;
            16'd6573: data <= 8'hF8;
            16'd6574: data <= 8'h00;
            16'd6575: data <= 8'hF8;
            16'd6576: data <= 8'h00;
            16'd6577: data <= 8'hF8;
            16'd6578: data <= 8'h00;
            16'd6579: data <= 8'hF8;
            16'd6580: data <= 8'h00;
            16'd6581: data <= 8'hF8;
            16'd6582: data <= 8'h00;
            16'd6583: data <= 8'hF8;
            16'd6584: data <= 8'h00;
            16'd6585: data <= 8'hF8;
            16'd6586: data <= 8'h00;
            16'd6587: data <= 8'hF8;
            16'd6588: data <= 8'h00;
            16'd6589: data <= 8'hF8;
            16'd6590: data <= 8'h00;
            16'd6591: data <= 8'hF8;
            16'd6592: data <= 8'h00;
            16'd6593: data <= 8'hF8;
            16'd6594: data <= 8'h00;
            16'd6595: data <= 8'hF8;
            16'd6596: data <= 8'h00;
            16'd6597: data <= 8'hF8;
            16'd6598: data <= 8'h00;
            16'd6599: data <= 8'hF8;
            16'd6600: data <= 8'hFF;
            16'd6601: data <= 8'hFF;
            16'd6602: data <= 8'h00;
            16'd6603: data <= 8'hF8;
            16'd6604: data <= 8'h00;
            16'd6605: data <= 8'hF8;
            16'd6606: data <= 8'h00;
            16'd6607: data <= 8'hF8;
            16'd6608: data <= 8'h00;
            16'd6609: data <= 8'hF8;
            16'd6610: data <= 8'h00;
            16'd6611: data <= 8'hF8;
            16'd6612: data <= 8'h00;
            16'd6613: data <= 8'hF8;
            16'd6614: data <= 8'h00;
            16'd6615: data <= 8'hF8;
            16'd6616: data <= 8'h00;
            16'd6617: data <= 8'hF8;
            16'd6618: data <= 8'h00;
            16'd6619: data <= 8'hF8;
            16'd6620: data <= 8'h00;
            16'd6621: data <= 8'hF8;
            16'd6622: data <= 8'h00;
            16'd6623: data <= 8'hF8;
            16'd6624: data <= 8'h00;
            16'd6625: data <= 8'hF8;
            16'd6626: data <= 8'h00;
            16'd6627: data <= 8'hF8;
            16'd6628: data <= 8'h00;
            16'd6629: data <= 8'hF8;
            16'd6630: data <= 8'h00;
            16'd6631: data <= 8'hF8;
            16'd6632: data <= 8'h00;
            16'd6633: data <= 8'hF8;
            16'd6634: data <= 8'h00;
            16'd6635: data <= 8'hF8;
            16'd6636: data <= 8'h00;
            16'd6637: data <= 8'hF8;
            16'd6638: data <= 8'h00;
            16'd6639: data <= 8'hF8;
            16'd6640: data <= 8'hFF;
            16'd6641: data <= 8'hFF;
            16'd6642: data <= 8'h00;
            16'd6643: data <= 8'hF8;
            16'd6644: data <= 8'h00;
            16'd6645: data <= 8'hF8;
            16'd6646: data <= 8'h00;
            16'd6647: data <= 8'hF8;
            16'd6648: data <= 8'h00;
            16'd6649: data <= 8'hF8;
            16'd6650: data <= 8'h00;
            16'd6651: data <= 8'hF8;
            16'd6652: data <= 8'h00;
            16'd6653: data <= 8'hF8;
            16'd6654: data <= 8'h00;
            16'd6655: data <= 8'hF8;
            16'd6656: data <= 8'h00;
            16'd6657: data <= 8'hF8;
            16'd6658: data <= 8'h00;
            16'd6659: data <= 8'hF8;
            16'd6660: data <= 8'h00;
            16'd6661: data <= 8'hF8;
            16'd6662: data <= 8'h00;
            16'd6663: data <= 8'hF8;
            16'd6664: data <= 8'h00;
            16'd6665: data <= 8'hF8;
            16'd6666: data <= 8'h00;
            16'd6667: data <= 8'hF8;
            16'd6668: data <= 8'h00;
            16'd6669: data <= 8'hF8;
            16'd6670: data <= 8'h00;
            16'd6671: data <= 8'hF8;
            16'd6672: data <= 8'h00;
            16'd6673: data <= 8'hF8;
            16'd6674: data <= 8'h00;
            16'd6675: data <= 8'hF8;
            16'd6676: data <= 8'h00;
            16'd6677: data <= 8'hF8;
            16'd6678: data <= 8'h00;
            16'd6679: data <= 8'hF8;
            16'd6680: data <= 8'hFF;
            16'd6681: data <= 8'hFF;
            16'd6682: data <= 8'h00;
            16'd6683: data <= 8'hF8;
            16'd6684: data <= 8'h00;
            16'd6685: data <= 8'hF8;
            16'd6686: data <= 8'h00;
            16'd6687: data <= 8'hF8;
            16'd6688: data <= 8'h00;
            16'd6689: data <= 8'hF8;
            16'd6690: data <= 8'h00;
            16'd6691: data <= 8'hF8;
            16'd6692: data <= 8'h00;
            16'd6693: data <= 8'hF8;
            16'd6694: data <= 8'h00;
            16'd6695: data <= 8'hF8;
            16'd6696: data <= 8'h00;
            16'd6697: data <= 8'hF8;
            16'd6698: data <= 8'h00;
            16'd6699: data <= 8'hF8;
            16'd6700: data <= 8'h00;
            16'd6701: data <= 8'hF8;
            16'd6702: data <= 8'h00;
            16'd6703: data <= 8'hF8;
            16'd6704: data <= 8'h00;
            16'd6705: data <= 8'hF8;
            16'd6706: data <= 8'h00;
            16'd6707: data <= 8'hF8;
            16'd6708: data <= 8'h00;
            16'd6709: data <= 8'hF8;
            16'd6710: data <= 8'h00;
            16'd6711: data <= 8'hF8;
            16'd6712: data <= 8'h00;
            16'd6713: data <= 8'hF8;
            16'd6714: data <= 8'h00;
            16'd6715: data <= 8'hF8;
            16'd6716: data <= 8'h00;
            16'd6717: data <= 8'hF8;
            16'd6718: data <= 8'h00;
            16'd6719: data <= 8'hF8;
            16'd6720: data <= 8'hFF;
            16'd6721: data <= 8'hFF;
            16'd6722: data <= 8'h00;
            16'd6723: data <= 8'hF8;
            16'd6724: data <= 8'h00;
            16'd6725: data <= 8'hF8;
            16'd6726: data <= 8'h00;
            16'd6727: data <= 8'hF8;
            16'd6728: data <= 8'h00;
            16'd6729: data <= 8'hF8;
            16'd6730: data <= 8'h00;
            16'd6731: data <= 8'hF8;
            16'd6732: data <= 8'h00;
            16'd6733: data <= 8'hF8;
            16'd6734: data <= 8'h00;
            16'd6735: data <= 8'hF8;
            16'd6736: data <= 8'h00;
            16'd6737: data <= 8'hF8;
            16'd6738: data <= 8'h00;
            16'd6739: data <= 8'hF8;
            16'd6740: data <= 8'h00;
            16'd6741: data <= 8'hF8;
            16'd6742: data <= 8'h00;
            16'd6743: data <= 8'hF8;
            16'd6744: data <= 8'h00;
            16'd6745: data <= 8'hF8;
            16'd6746: data <= 8'h00;
            16'd6747: data <= 8'hF8;
            16'd6748: data <= 8'h00;
            16'd6749: data <= 8'hF8;
            16'd6750: data <= 8'h00;
            16'd6751: data <= 8'hF8;
            16'd6752: data <= 8'h00;
            16'd6753: data <= 8'hF8;
            16'd6754: data <= 8'h00;
            16'd6755: data <= 8'hF8;
            16'd6756: data <= 8'h00;
            16'd6757: data <= 8'hF8;
            16'd6758: data <= 8'h00;
            16'd6759: data <= 8'hF8;
            16'd6760: data <= 8'hFF;
            16'd6761: data <= 8'hFF;
            16'd6762: data <= 8'h00;
            16'd6763: data <= 8'hF8;
            16'd6764: data <= 8'h00;
            16'd6765: data <= 8'hF8;
            16'd6766: data <= 8'h00;
            16'd6767: data <= 8'hF8;
            16'd6768: data <= 8'h00;
            16'd6769: data <= 8'hF8;
            16'd6770: data <= 8'h00;
            16'd6771: data <= 8'hF8;
            16'd6772: data <= 8'h00;
            16'd6773: data <= 8'hF8;
            16'd6774: data <= 8'h00;
            16'd6775: data <= 8'hF8;
            16'd6776: data <= 8'h00;
            16'd6777: data <= 8'hF8;
            16'd6778: data <= 8'h00;
            16'd6779: data <= 8'hF8;
            16'd6780: data <= 8'h00;
            16'd6781: data <= 8'hF8;
            16'd6782: data <= 8'h00;
            16'd6783: data <= 8'hF8;
            16'd6784: data <= 8'h00;
            16'd6785: data <= 8'hF8;
            16'd6786: data <= 8'h00;
            16'd6787: data <= 8'hF8;
            16'd6788: data <= 8'h00;
            16'd6789: data <= 8'hF8;
            16'd6790: data <= 8'h00;
            16'd6791: data <= 8'hF8;
            16'd6792: data <= 8'h00;
            16'd6793: data <= 8'hF8;
            16'd6794: data <= 8'h00;
            16'd6795: data <= 8'hF8;
            16'd6796: data <= 8'h00;
            16'd6797: data <= 8'hF8;
            16'd6798: data <= 8'h00;
            16'd6799: data <= 8'hF8;
            16'd6800: data <= 8'hFF;
            16'd6801: data <= 8'hFF;
            16'd6802: data <= 8'h00;
            16'd6803: data <= 8'hF8;
            16'd6804: data <= 8'h00;
            16'd6805: data <= 8'hF8;
            16'd6806: data <= 8'h00;
            16'd6807: data <= 8'hF8;
            16'd6808: data <= 8'h00;
            16'd6809: data <= 8'hF8;
            16'd6810: data <= 8'h00;
            16'd6811: data <= 8'hF8;
            16'd6812: data <= 8'h00;
            16'd6813: data <= 8'hF8;
            16'd6814: data <= 8'h00;
            16'd6815: data <= 8'hF8;
            16'd6816: data <= 8'h00;
            16'd6817: data <= 8'hF8;
            16'd6818: data <= 8'h00;
            16'd6819: data <= 8'hF8;
            16'd6820: data <= 8'h00;
            16'd6821: data <= 8'hF8;
            16'd6822: data <= 8'h00;
            16'd6823: data <= 8'hF8;
            16'd6824: data <= 8'h00;
            16'd6825: data <= 8'hF8;
            16'd6826: data <= 8'h00;
            16'd6827: data <= 8'hF8;
            16'd6828: data <= 8'h00;
            16'd6829: data <= 8'hF8;
            16'd6830: data <= 8'h00;
            16'd6831: data <= 8'hF8;
            16'd6832: data <= 8'h00;
            16'd6833: data <= 8'hF8;
            16'd6834: data <= 8'h00;
            16'd6835: data <= 8'hF8;
            16'd6836: data <= 8'h00;
            16'd6837: data <= 8'hF8;
            16'd6838: data <= 8'h00;
            16'd6839: data <= 8'hF8;
            16'd6840: data <= 8'hFF;
            16'd6841: data <= 8'hFF;
            16'd6842: data <= 8'h00;
            16'd6843: data <= 8'hF8;
            16'd6844: data <= 8'h00;
            16'd6845: data <= 8'hF8;
            16'd6846: data <= 8'h00;
            16'd6847: data <= 8'hF8;
            16'd6848: data <= 8'h00;
            16'd6849: data <= 8'hF8;
            16'd6850: data <= 8'h00;
            16'd6851: data <= 8'hF8;
            16'd6852: data <= 8'h00;
            16'd6853: data <= 8'hF8;
            16'd6854: data <= 8'h00;
            16'd6855: data <= 8'hF8;
            16'd6856: data <= 8'h00;
            16'd6857: data <= 8'hF8;
            16'd6858: data <= 8'h00;
            16'd6859: data <= 8'hF8;
            16'd6860: data <= 8'h00;
            16'd6861: data <= 8'hF8;
            16'd6862: data <= 8'h00;
            16'd6863: data <= 8'hF8;
            16'd6864: data <= 8'h00;
            16'd6865: data <= 8'hF8;
            16'd6866: data <= 8'h00;
            16'd6867: data <= 8'hF8;
            16'd6868: data <= 8'h00;
            16'd6869: data <= 8'hF8;
            16'd6870: data <= 8'h00;
            16'd6871: data <= 8'hF8;
            16'd6872: data <= 8'h00;
            16'd6873: data <= 8'hF8;
            16'd6874: data <= 8'h00;
            16'd6875: data <= 8'hF8;
            16'd6876: data <= 8'h00;
            16'd6877: data <= 8'hF8;
            16'd6878: data <= 8'h00;
            16'd6879: data <= 8'hF8;
            16'd6880: data <= 8'hFF;
            16'd6881: data <= 8'hFF;
            16'd6882: data <= 8'h00;
            16'd6883: data <= 8'hF8;
            16'd6884: data <= 8'h00;
            16'd6885: data <= 8'hF8;
            16'd6886: data <= 8'h00;
            16'd6887: data <= 8'hF8;
            16'd6888: data <= 8'h00;
            16'd6889: data <= 8'hF8;
            16'd6890: data <= 8'h00;
            16'd6891: data <= 8'hF8;
            16'd6892: data <= 8'h00;
            16'd6893: data <= 8'hF8;
            16'd6894: data <= 8'h00;
            16'd6895: data <= 8'hF8;
            16'd6896: data <= 8'h00;
            16'd6897: data <= 8'hF8;
            16'd6898: data <= 8'h00;
            16'd6899: data <= 8'hF8;
            16'd6900: data <= 8'h00;
            16'd6901: data <= 8'hF8;
            16'd6902: data <= 8'h00;
            16'd6903: data <= 8'hF8;
            16'd6904: data <= 8'h00;
            16'd6905: data <= 8'hF8;
            16'd6906: data <= 8'h00;
            16'd6907: data <= 8'hF8;
            16'd6908: data <= 8'h00;
            16'd6909: data <= 8'hF8;
            16'd6910: data <= 8'h00;
            16'd6911: data <= 8'hF8;
            16'd6912: data <= 8'h00;
            16'd6913: data <= 8'hF8;
            16'd6914: data <= 8'h00;
            16'd6915: data <= 8'hF8;
            16'd6916: data <= 8'h00;
            16'd6917: data <= 8'hF8;
            16'd6918: data <= 8'h00;
            16'd6919: data <= 8'hF8;
            16'd6920: data <= 8'hFF;
            16'd6921: data <= 8'hFF;
            16'd6922: data <= 8'h00;
            16'd6923: data <= 8'hF8;
            16'd6924: data <= 8'h00;
            16'd6925: data <= 8'hF8;
            16'd6926: data <= 8'h00;
            16'd6927: data <= 8'hF8;
            16'd6928: data <= 8'h00;
            16'd6929: data <= 8'hF8;
            16'd6930: data <= 8'h00;
            16'd6931: data <= 8'hF8;
            16'd6932: data <= 8'h00;
            16'd6933: data <= 8'hF8;
            16'd6934: data <= 8'h00;
            16'd6935: data <= 8'hF8;
            16'd6936: data <= 8'h00;
            16'd6937: data <= 8'hF8;
            16'd6938: data <= 8'h00;
            16'd6939: data <= 8'hF8;
            16'd6940: data <= 8'h00;
            16'd6941: data <= 8'hF8;
            16'd6942: data <= 8'h00;
            16'd6943: data <= 8'hF8;
            16'd6944: data <= 8'h00;
            16'd6945: data <= 8'hF8;
            16'd6946: data <= 8'h00;
            16'd6947: data <= 8'hF8;
            16'd6948: data <= 8'h00;
            16'd6949: data <= 8'hF8;
            16'd6950: data <= 8'h00;
            16'd6951: data <= 8'hF8;
            16'd6952: data <= 8'h00;
            16'd6953: data <= 8'hF8;
            16'd6954: data <= 8'h00;
            16'd6955: data <= 8'hF8;
            16'd6956: data <= 8'h00;
            16'd6957: data <= 8'hF8;
            16'd6958: data <= 8'h00;
            16'd6959: data <= 8'hF8;
            16'd6960: data <= 8'hFF;
            16'd6961: data <= 8'hFF;
            16'd6962: data <= 8'h00;
            16'd6963: data <= 8'hF8;
            16'd6964: data <= 8'h00;
            16'd6965: data <= 8'hF8;
            16'd6966: data <= 8'h00;
            16'd6967: data <= 8'hF8;
            16'd6968: data <= 8'h00;
            16'd6969: data <= 8'hF8;
            16'd6970: data <= 8'h00;
            16'd6971: data <= 8'hF8;
            16'd6972: data <= 8'h00;
            16'd6973: data <= 8'hF8;
            16'd6974: data <= 8'h00;
            16'd6975: data <= 8'hF8;
            16'd6976: data <= 8'h00;
            16'd6977: data <= 8'hF8;
            16'd6978: data <= 8'h00;
            16'd6979: data <= 8'hF8;
            16'd6980: data <= 8'h00;
            16'd6981: data <= 8'hF8;
            16'd6982: data <= 8'h00;
            16'd6983: data <= 8'hF8;
            16'd6984: data <= 8'h00;
            16'd6985: data <= 8'hF8;
            16'd6986: data <= 8'h00;
            16'd6987: data <= 8'hF8;
            16'd6988: data <= 8'h00;
            16'd6989: data <= 8'hF8;
            16'd6990: data <= 8'h00;
            16'd6991: data <= 8'hF8;
            16'd6992: data <= 8'h00;
            16'd6993: data <= 8'hF8;
            16'd6994: data <= 8'h00;
            16'd6995: data <= 8'hF8;
            16'd6996: data <= 8'h00;
            16'd6997: data <= 8'hF8;
            16'd6998: data <= 8'h00;
            16'd6999: data <= 8'hF8;
            16'd7000: data <= 8'hFF;
            16'd7001: data <= 8'hFF;
            16'd7002: data <= 8'h00;
            16'd7003: data <= 8'hF8;
            16'd7004: data <= 8'h00;
            16'd7005: data <= 8'hF8;
            16'd7006: data <= 8'h00;
            16'd7007: data <= 8'hF8;
            16'd7008: data <= 8'h00;
            16'd7009: data <= 8'hF8;
            16'd7010: data <= 8'h00;
            16'd7011: data <= 8'hF8;
            16'd7012: data <= 8'h00;
            16'd7013: data <= 8'hF8;
            16'd7014: data <= 8'h00;
            16'd7015: data <= 8'hF8;
            16'd7016: data <= 8'h00;
            16'd7017: data <= 8'hF8;
            16'd7018: data <= 8'h00;
            16'd7019: data <= 8'hF8;
            16'd7020: data <= 8'h00;
            16'd7021: data <= 8'hF8;
            16'd7022: data <= 8'h00;
            16'd7023: data <= 8'hF8;
            16'd7024: data <= 8'h00;
            16'd7025: data <= 8'hF8;
            16'd7026: data <= 8'h00;
            16'd7027: data <= 8'hF8;
            16'd7028: data <= 8'h00;
            16'd7029: data <= 8'hF8;
            16'd7030: data <= 8'h00;
            16'd7031: data <= 8'hF8;
            16'd7032: data <= 8'h00;
            16'd7033: data <= 8'hF8;
            16'd7034: data <= 8'h00;
            16'd7035: data <= 8'hF8;
            16'd7036: data <= 8'h00;
            16'd7037: data <= 8'hF8;
            16'd7038: data <= 8'h00;
            16'd7039: data <= 8'hF8;
            16'd7040: data <= 8'hFF;
            16'd7041: data <= 8'hFF;
            16'd7042: data <= 8'h00;
            16'd7043: data <= 8'hF8;
            16'd7044: data <= 8'h00;
            16'd7045: data <= 8'hF8;
            16'd7046: data <= 8'h00;
            16'd7047: data <= 8'hF8;
            16'd7048: data <= 8'h00;
            16'd7049: data <= 8'hF8;
            16'd7050: data <= 8'h00;
            16'd7051: data <= 8'hF8;
            16'd7052: data <= 8'h00;
            16'd7053: data <= 8'hF8;
            16'd7054: data <= 8'h00;
            16'd7055: data <= 8'hF8;
            16'd7056: data <= 8'h00;
            16'd7057: data <= 8'hF8;
            16'd7058: data <= 8'h00;
            16'd7059: data <= 8'hF8;
            16'd7060: data <= 8'h00;
            16'd7061: data <= 8'hF8;
            16'd7062: data <= 8'h00;
            16'd7063: data <= 8'hF8;
            16'd7064: data <= 8'h00;
            16'd7065: data <= 8'hF8;
            16'd7066: data <= 8'h00;
            16'd7067: data <= 8'hF8;
            16'd7068: data <= 8'h00;
            16'd7069: data <= 8'hF8;
            16'd7070: data <= 8'h00;
            16'd7071: data <= 8'hF8;
            16'd7072: data <= 8'h00;
            16'd7073: data <= 8'hF8;
            16'd7074: data <= 8'h00;
            16'd7075: data <= 8'hF8;
            16'd7076: data <= 8'h00;
            16'd7077: data <= 8'hF8;
            16'd7078: data <= 8'h00;
            16'd7079: data <= 8'hF8;
            16'd7080: data <= 8'hFF;
            16'd7081: data <= 8'hFF;
            16'd7082: data <= 8'h00;
            16'd7083: data <= 8'hF8;
            16'd7084: data <= 8'h00;
            16'd7085: data <= 8'hF8;
            16'd7086: data <= 8'h00;
            16'd7087: data <= 8'hF8;
            16'd7088: data <= 8'h00;
            16'd7089: data <= 8'hF8;
            16'd7090: data <= 8'h00;
            16'd7091: data <= 8'hF8;
            16'd7092: data <= 8'h00;
            16'd7093: data <= 8'hF8;
            16'd7094: data <= 8'h00;
            16'd7095: data <= 8'hF8;
            16'd7096: data <= 8'h00;
            16'd7097: data <= 8'hF8;
            16'd7098: data <= 8'h00;
            16'd7099: data <= 8'hF8;
            16'd7100: data <= 8'h00;
            16'd7101: data <= 8'hF8;
            16'd7102: data <= 8'h00;
            16'd7103: data <= 8'hF8;
            16'd7104: data <= 8'h00;
            16'd7105: data <= 8'hF8;
            16'd7106: data <= 8'h00;
            16'd7107: data <= 8'hF8;
            16'd7108: data <= 8'h00;
            16'd7109: data <= 8'hF8;
            16'd7110: data <= 8'h00;
            16'd7111: data <= 8'hF8;
            16'd7112: data <= 8'h00;
            16'd7113: data <= 8'hF8;
            16'd7114: data <= 8'h00;
            16'd7115: data <= 8'hF8;
            16'd7116: data <= 8'h00;
            16'd7117: data <= 8'hF8;
            16'd7118: data <= 8'h00;
            16'd7119: data <= 8'hF8;
            16'd7120: data <= 8'hFF;
            16'd7121: data <= 8'hFF;
            16'd7122: data <= 8'h00;
            16'd7123: data <= 8'hF8;
            16'd7124: data <= 8'h00;
            16'd7125: data <= 8'hF8;
            16'd7126: data <= 8'h00;
            16'd7127: data <= 8'hF8;
            16'd7128: data <= 8'h00;
            16'd7129: data <= 8'hF8;
            16'd7130: data <= 8'h00;
            16'd7131: data <= 8'hF8;
            16'd7132: data <= 8'h00;
            16'd7133: data <= 8'hF8;
            16'd7134: data <= 8'h00;
            16'd7135: data <= 8'hF8;
            16'd7136: data <= 8'h00;
            16'd7137: data <= 8'hF8;
            16'd7138: data <= 8'h00;
            16'd7139: data <= 8'hF8;
            16'd7140: data <= 8'h00;
            16'd7141: data <= 8'hF8;
            16'd7142: data <= 8'h00;
            16'd7143: data <= 8'hF8;
            16'd7144: data <= 8'h00;
            16'd7145: data <= 8'hF8;
            16'd7146: data <= 8'h00;
            16'd7147: data <= 8'hF8;
            16'd7148: data <= 8'h00;
            16'd7149: data <= 8'hF8;
            16'd7150: data <= 8'h00;
            16'd7151: data <= 8'hF8;
            16'd7152: data <= 8'h00;
            16'd7153: data <= 8'hF8;
            16'd7154: data <= 8'h00;
            16'd7155: data <= 8'hF8;
            16'd7156: data <= 8'h00;
            16'd7157: data <= 8'hF8;
            16'd7158: data <= 8'h00;
            16'd7159: data <= 8'hF8;
            16'd7160: data <= 8'hFF;
            16'd7161: data <= 8'hFF;
            16'd7162: data <= 8'h00;
            16'd7163: data <= 8'hF8;
            16'd7164: data <= 8'h00;
            16'd7165: data <= 8'hF8;
            16'd7166: data <= 8'h00;
            16'd7167: data <= 8'hF8;
            16'd7168: data <= 8'h00;
            16'd7169: data <= 8'hF8;
            16'd7170: data <= 8'h00;
            16'd7171: data <= 8'hF8;
            16'd7172: data <= 8'h00;
            16'd7173: data <= 8'hF8;
            16'd7174: data <= 8'h00;
            16'd7175: data <= 8'hF8;
            16'd7176: data <= 8'h00;
            16'd7177: data <= 8'hF8;
            16'd7178: data <= 8'h00;
            16'd7179: data <= 8'hF8;
            16'd7180: data <= 8'h00;
            16'd7181: data <= 8'hF8;
            16'd7182: data <= 8'h00;
            16'd7183: data <= 8'hF8;
            16'd7184: data <= 8'h00;
            16'd7185: data <= 8'hF8;
            16'd7186: data <= 8'h00;
            16'd7187: data <= 8'hF8;
            16'd7188: data <= 8'h00;
            16'd7189: data <= 8'hF8;
            16'd7190: data <= 8'h00;
            16'd7191: data <= 8'hF8;
            16'd7192: data <= 8'h00;
            16'd7193: data <= 8'hF8;
            16'd7194: data <= 8'h00;
            16'd7195: data <= 8'hF8;
            16'd7196: data <= 8'h00;
            16'd7197: data <= 8'hF8;
            16'd7198: data <= 8'h00;
            16'd7199: data <= 8'hF8;
            16'd7200: data <= 8'hFF;
            16'd7201: data <= 8'hFF;
            16'd7202: data <= 8'h00;
            16'd7203: data <= 8'hF8;
            16'd7204: data <= 8'h00;
            16'd7205: data <= 8'hF8;
            16'd7206: data <= 8'h00;
            16'd7207: data <= 8'hF8;
            16'd7208: data <= 8'h00;
            16'd7209: data <= 8'hF8;
            16'd7210: data <= 8'h00;
            16'd7211: data <= 8'hF8;
            16'd7212: data <= 8'h00;
            16'd7213: data <= 8'hF8;
            16'd7214: data <= 8'h00;
            16'd7215: data <= 8'hF8;
            16'd7216: data <= 8'h00;
            16'd7217: data <= 8'hF8;
            16'd7218: data <= 8'h00;
            16'd7219: data <= 8'hF8;
            16'd7220: data <= 8'h00;
            16'd7221: data <= 8'hF8;
            16'd7222: data <= 8'h00;
            16'd7223: data <= 8'hF8;
            16'd7224: data <= 8'h00;
            16'd7225: data <= 8'hF8;
            16'd7226: data <= 8'h00;
            16'd7227: data <= 8'hF8;
            16'd7228: data <= 8'h00;
            16'd7229: data <= 8'hF8;
            16'd7230: data <= 8'h00;
            16'd7231: data <= 8'hF8;
            16'd7232: data <= 8'h00;
            16'd7233: data <= 8'hF8;
            16'd7234: data <= 8'h00;
            16'd7235: data <= 8'hF8;
            16'd7236: data <= 8'h00;
            16'd7237: data <= 8'hF8;
            16'd7238: data <= 8'h00;
            16'd7239: data <= 8'hF8;
            16'd7240: data <= 8'hFF;
            16'd7241: data <= 8'hFF;
            16'd7242: data <= 8'h00;
            16'd7243: data <= 8'hF8;
            16'd7244: data <= 8'h00;
            16'd7245: data <= 8'hF8;
            16'd7246: data <= 8'h00;
            16'd7247: data <= 8'hF8;
            16'd7248: data <= 8'h00;
            16'd7249: data <= 8'hF8;
            16'd7250: data <= 8'h00;
            16'd7251: data <= 8'hF8;
            16'd7252: data <= 8'h00;
            16'd7253: data <= 8'hF8;
            16'd7254: data <= 8'h00;
            16'd7255: data <= 8'hF8;
            16'd7256: data <= 8'h00;
            16'd7257: data <= 8'hF8;
            16'd7258: data <= 8'h00;
            16'd7259: data <= 8'hF8;
            16'd7260: data <= 8'h00;
            16'd7261: data <= 8'hF8;
            16'd7262: data <= 8'h00;
            16'd7263: data <= 8'hF8;
            16'd7264: data <= 8'h00;
            16'd7265: data <= 8'hF8;
            16'd7266: data <= 8'h00;
            16'd7267: data <= 8'hF8;
            16'd7268: data <= 8'h00;
            16'd7269: data <= 8'hF8;
            16'd7270: data <= 8'h00;
            16'd7271: data <= 8'hF8;
            16'd7272: data <= 8'h00;
            16'd7273: data <= 8'hF8;
            16'd7274: data <= 8'h00;
            16'd7275: data <= 8'hF8;
            16'd7276: data <= 8'h00;
            16'd7277: data <= 8'hF8;
            16'd7278: data <= 8'h00;
            16'd7279: data <= 8'hF8;
            16'd7280: data <= 8'hFF;
            16'd7281: data <= 8'hFF;
            16'd7282: data <= 8'h00;
            16'd7283: data <= 8'hF8;
            16'd7284: data <= 8'h00;
            16'd7285: data <= 8'hF8;
            16'd7286: data <= 8'h00;
            16'd7287: data <= 8'hF8;
            16'd7288: data <= 8'h00;
            16'd7289: data <= 8'hF8;
            16'd7290: data <= 8'h00;
            16'd7291: data <= 8'hF8;
            16'd7292: data <= 8'h00;
            16'd7293: data <= 8'hF8;
            16'd7294: data <= 8'h00;
            16'd7295: data <= 8'hF8;
            16'd7296: data <= 8'h00;
            16'd7297: data <= 8'hF8;
            16'd7298: data <= 8'h00;
            16'd7299: data <= 8'hF8;
            16'd7300: data <= 8'h00;
            16'd7301: data <= 8'hF8;
            16'd7302: data <= 8'h00;
            16'd7303: data <= 8'hF8;
            16'd7304: data <= 8'h00;
            16'd7305: data <= 8'hF8;
            16'd7306: data <= 8'h00;
            16'd7307: data <= 8'hF8;
            16'd7308: data <= 8'h00;
            16'd7309: data <= 8'hF8;
            16'd7310: data <= 8'h00;
            16'd7311: data <= 8'hF8;
            16'd7312: data <= 8'h00;
            16'd7313: data <= 8'hF8;
            16'd7314: data <= 8'h00;
            16'd7315: data <= 8'hF8;
            16'd7316: data <= 8'h00;
            16'd7317: data <= 8'hF8;
            16'd7318: data <= 8'h00;
            16'd7319: data <= 8'hF8;
            16'd7320: data <= 8'hFF;
            16'd7321: data <= 8'hFF;
            16'd7322: data <= 8'h00;
            16'd7323: data <= 8'hF8;
            16'd7324: data <= 8'h00;
            16'd7325: data <= 8'hF8;
            16'd7326: data <= 8'h00;
            16'd7327: data <= 8'hF8;
            16'd7328: data <= 8'h00;
            16'd7329: data <= 8'hF8;
            16'd7330: data <= 8'h00;
            16'd7331: data <= 8'hF8;
            16'd7332: data <= 8'h00;
            16'd7333: data <= 8'hF8;
            16'd7334: data <= 8'h00;
            16'd7335: data <= 8'hF8;
            16'd7336: data <= 8'h00;
            16'd7337: data <= 8'hF8;
            16'd7338: data <= 8'h00;
            16'd7339: data <= 8'hF8;
            16'd7340: data <= 8'h00;
            16'd7341: data <= 8'hF8;
            16'd7342: data <= 8'h00;
            16'd7343: data <= 8'hF8;
            16'd7344: data <= 8'h00;
            16'd7345: data <= 8'hF8;
            16'd7346: data <= 8'h00;
            16'd7347: data <= 8'hF8;
            16'd7348: data <= 8'h00;
            16'd7349: data <= 8'hF8;
            16'd7350: data <= 8'h00;
            16'd7351: data <= 8'hF8;
            16'd7352: data <= 8'h00;
            16'd7353: data <= 8'hF8;
            16'd7354: data <= 8'h00;
            16'd7355: data <= 8'hF8;
            16'd7356: data <= 8'h00;
            16'd7357: data <= 8'hF8;
            16'd7358: data <= 8'h00;
            16'd7359: data <= 8'hF8;
            16'd7360: data <= 8'hFF;
            16'd7361: data <= 8'hFF;
            16'd7362: data <= 8'h00;
            16'd7363: data <= 8'hF8;
            16'd7364: data <= 8'h00;
            16'd7365: data <= 8'hF8;
            16'd7366: data <= 8'h00;
            16'd7367: data <= 8'hF8;
            16'd7368: data <= 8'h00;
            16'd7369: data <= 8'hF8;
            16'd7370: data <= 8'h00;
            16'd7371: data <= 8'hF8;
            16'd7372: data <= 8'h00;
            16'd7373: data <= 8'hF8;
            16'd7374: data <= 8'h00;
            16'd7375: data <= 8'hF8;
            16'd7376: data <= 8'h00;
            16'd7377: data <= 8'hF8;
            16'd7378: data <= 8'h00;
            16'd7379: data <= 8'hF8;
            16'd7380: data <= 8'h00;
            16'd7381: data <= 8'hF8;
            16'd7382: data <= 8'h00;
            16'd7383: data <= 8'hF8;
            16'd7384: data <= 8'h00;
            16'd7385: data <= 8'hF8;
            16'd7386: data <= 8'h00;
            16'd7387: data <= 8'hF8;
            16'd7388: data <= 8'h00;
            16'd7389: data <= 8'hF8;
            16'd7390: data <= 8'h00;
            16'd7391: data <= 8'hF8;
            16'd7392: data <= 8'h00;
            16'd7393: data <= 8'hF8;
            16'd7394: data <= 8'h00;
            16'd7395: data <= 8'hF8;
            16'd7396: data <= 8'h00;
            16'd7397: data <= 8'hF8;
            16'd7398: data <= 8'h00;
            16'd7399: data <= 8'hF8;
            16'd7400: data <= 8'hFF;
            16'd7401: data <= 8'hFF;
            16'd7402: data <= 8'h00;
            16'd7403: data <= 8'hF8;
            16'd7404: data <= 8'h00;
            16'd7405: data <= 8'hF8;
            16'd7406: data <= 8'h00;
            16'd7407: data <= 8'hF8;
            16'd7408: data <= 8'h00;
            16'd7409: data <= 8'hF8;
            16'd7410: data <= 8'h00;
            16'd7411: data <= 8'hF8;
            16'd7412: data <= 8'h00;
            16'd7413: data <= 8'hF8;
            16'd7414: data <= 8'h00;
            16'd7415: data <= 8'hF8;
            16'd7416: data <= 8'h00;
            16'd7417: data <= 8'hF8;
            16'd7418: data <= 8'h00;
            16'd7419: data <= 8'hF8;
            16'd7420: data <= 8'h00;
            16'd7421: data <= 8'hF8;
            16'd7422: data <= 8'h00;
            16'd7423: data <= 8'hF8;
            16'd7424: data <= 8'h00;
            16'd7425: data <= 8'hF8;
            16'd7426: data <= 8'h00;
            16'd7427: data <= 8'hF8;
            16'd7428: data <= 8'h00;
            16'd7429: data <= 8'hF8;
            16'd7430: data <= 8'h00;
            16'd7431: data <= 8'hF8;
            16'd7432: data <= 8'h00;
            16'd7433: data <= 8'hF8;
            16'd7434: data <= 8'h00;
            16'd7435: data <= 8'hF8;
            16'd7436: data <= 8'h00;
            16'd7437: data <= 8'hF8;
            16'd7438: data <= 8'h00;
            16'd7439: data <= 8'hF8;
            16'd7440: data <= 8'hFF;
            16'd7441: data <= 8'hFF;
            16'd7442: data <= 8'h00;
            16'd7443: data <= 8'hF8;
            16'd7444: data <= 8'h00;
            16'd7445: data <= 8'hF8;
            16'd7446: data <= 8'h00;
            16'd7447: data <= 8'hF8;
            16'd7448: data <= 8'h00;
            16'd7449: data <= 8'hF8;
            16'd7450: data <= 8'h00;
            16'd7451: data <= 8'hF8;
            16'd7452: data <= 8'h00;
            16'd7453: data <= 8'hF8;
            16'd7454: data <= 8'h00;
            16'd7455: data <= 8'hF8;
            16'd7456: data <= 8'h00;
            16'd7457: data <= 8'hF8;
            16'd7458: data <= 8'h00;
            16'd7459: data <= 8'hF8;
            16'd7460: data <= 8'h00;
            16'd7461: data <= 8'hF8;
            16'd7462: data <= 8'h00;
            16'd7463: data <= 8'hF8;
            16'd7464: data <= 8'h00;
            16'd7465: data <= 8'hF8;
            16'd7466: data <= 8'h00;
            16'd7467: data <= 8'hF8;
            16'd7468: data <= 8'h00;
            16'd7469: data <= 8'hF8;
            16'd7470: data <= 8'h00;
            16'd7471: data <= 8'hF8;
            16'd7472: data <= 8'h00;
            16'd7473: data <= 8'hF8;
            16'd7474: data <= 8'h00;
            16'd7475: data <= 8'hF8;
            16'd7476: data <= 8'h00;
            16'd7477: data <= 8'hF8;
            16'd7478: data <= 8'h00;
            16'd7479: data <= 8'hF8;
            16'd7480: data <= 8'hFF;
            16'd7481: data <= 8'hFF;
            16'd7482: data <= 8'h00;
            16'd7483: data <= 8'hF8;
            16'd7484: data <= 8'h00;
            16'd7485: data <= 8'hF8;
            16'd7486: data <= 8'h00;
            16'd7487: data <= 8'hF8;
            16'd7488: data <= 8'h00;
            16'd7489: data <= 8'hF8;
            16'd7490: data <= 8'h00;
            16'd7491: data <= 8'hF8;
            16'd7492: data <= 8'h00;
            16'd7493: data <= 8'hF8;
            16'd7494: data <= 8'h00;
            16'd7495: data <= 8'hF8;
            16'd7496: data <= 8'h00;
            16'd7497: data <= 8'hF8;
            16'd7498: data <= 8'h00;
            16'd7499: data <= 8'hF8;
            16'd7500: data <= 8'h00;
            16'd7501: data <= 8'hF8;
            16'd7502: data <= 8'h00;
            16'd7503: data <= 8'hF8;
            16'd7504: data <= 8'h00;
            16'd7505: data <= 8'hF8;
            16'd7506: data <= 8'h00;
            16'd7507: data <= 8'hF8;
            16'd7508: data <= 8'h00;
            16'd7509: data <= 8'hF8;
            16'd7510: data <= 8'h00;
            16'd7511: data <= 8'hF8;
            16'd7512: data <= 8'h00;
            16'd7513: data <= 8'hF8;
            16'd7514: data <= 8'h00;
            16'd7515: data <= 8'hF8;
            16'd7516: data <= 8'h00;
            16'd7517: data <= 8'hF8;
            16'd7518: data <= 8'h00;
            16'd7519: data <= 8'hF8;
            16'd7520: data <= 8'hFF;
            16'd7521: data <= 8'hFF;
            16'd7522: data <= 8'h00;
            16'd7523: data <= 8'hF8;
            16'd7524: data <= 8'h00;
            16'd7525: data <= 8'hF8;
            16'd7526: data <= 8'h00;
            16'd7527: data <= 8'hF8;
            16'd7528: data <= 8'h00;
            16'd7529: data <= 8'hF8;
            16'd7530: data <= 8'h00;
            16'd7531: data <= 8'hF8;
            16'd7532: data <= 8'h00;
            16'd7533: data <= 8'hF8;
            16'd7534: data <= 8'h00;
            16'd7535: data <= 8'hF8;
            16'd7536: data <= 8'h00;
            16'd7537: data <= 8'hF8;
            16'd7538: data <= 8'h00;
            16'd7539: data <= 8'hF8;
            16'd7540: data <= 8'h00;
            16'd7541: data <= 8'hF8;
            16'd7542: data <= 8'h00;
            16'd7543: data <= 8'hF8;
            16'd7544: data <= 8'h00;
            16'd7545: data <= 8'hF8;
            16'd7546: data <= 8'h00;
            16'd7547: data <= 8'hF8;
            16'd7548: data <= 8'h00;
            16'd7549: data <= 8'hF8;
            16'd7550: data <= 8'h00;
            16'd7551: data <= 8'hF8;
            16'd7552: data <= 8'h00;
            16'd7553: data <= 8'hF8;
            16'd7554: data <= 8'h00;
            16'd7555: data <= 8'hF8;
            16'd7556: data <= 8'h00;
            16'd7557: data <= 8'hF8;
            16'd7558: data <= 8'h00;
            16'd7559: data <= 8'hF8;
            16'd7560: data <= 8'hFF;
            16'd7561: data <= 8'hFF;
            16'd7562: data <= 8'h00;
            16'd7563: data <= 8'hF8;
            16'd7564: data <= 8'h00;
            16'd7565: data <= 8'hF8;
            16'd7566: data <= 8'h00;
            16'd7567: data <= 8'hF8;
            16'd7568: data <= 8'h00;
            16'd7569: data <= 8'hF8;
            16'd7570: data <= 8'h00;
            16'd7571: data <= 8'hF8;
            16'd7572: data <= 8'h00;
            16'd7573: data <= 8'hF8;
            16'd7574: data <= 8'h00;
            16'd7575: data <= 8'hF8;
            16'd7576: data <= 8'h00;
            16'd7577: data <= 8'hF8;
            16'd7578: data <= 8'h00;
            16'd7579: data <= 8'hF8;
            16'd7580: data <= 8'h00;
            16'd7581: data <= 8'hF8;
            16'd7582: data <= 8'h00;
            16'd7583: data <= 8'hF8;
            16'd7584: data <= 8'h00;
            16'd7585: data <= 8'hF8;
            16'd7586: data <= 8'h00;
            16'd7587: data <= 8'hF8;
            16'd7588: data <= 8'h00;
            16'd7589: data <= 8'hF8;
            16'd7590: data <= 8'h00;
            16'd7591: data <= 8'hF8;
            16'd7592: data <= 8'h00;
            16'd7593: data <= 8'hF8;
            16'd7594: data <= 8'h00;
            16'd7595: data <= 8'hF8;
            16'd7596: data <= 8'h00;
            16'd7597: data <= 8'hF8;
            16'd7598: data <= 8'h00;
            16'd7599: data <= 8'hF8;
            16'd7600: data <= 8'hFF;
            16'd7601: data <= 8'hFF;
            16'd7602: data <= 8'h00;
            16'd7603: data <= 8'hF8;
            16'd7604: data <= 8'h00;
            16'd7605: data <= 8'hF8;
            16'd7606: data <= 8'h00;
            16'd7607: data <= 8'hF8;
            16'd7608: data <= 8'h00;
            16'd7609: data <= 8'hF8;
            16'd7610: data <= 8'h00;
            16'd7611: data <= 8'hF8;
            16'd7612: data <= 8'h00;
            16'd7613: data <= 8'hF8;
            16'd7614: data <= 8'h00;
            16'd7615: data <= 8'hF8;
            16'd7616: data <= 8'h00;
            16'd7617: data <= 8'hF8;
            16'd7618: data <= 8'h00;
            16'd7619: data <= 8'hF8;
            16'd7620: data <= 8'h00;
            16'd7621: data <= 8'hF8;
            16'd7622: data <= 8'h00;
            16'd7623: data <= 8'hF8;
            16'd7624: data <= 8'h00;
            16'd7625: data <= 8'hF8;
            16'd7626: data <= 8'h00;
            16'd7627: data <= 8'hF8;
            16'd7628: data <= 8'h00;
            16'd7629: data <= 8'hF8;
            16'd7630: data <= 8'h00;
            16'd7631: data <= 8'hF8;
            16'd7632: data <= 8'h00;
            16'd7633: data <= 8'hF8;
            16'd7634: data <= 8'h00;
            16'd7635: data <= 8'hF8;
            16'd7636: data <= 8'h00;
            16'd7637: data <= 8'hF8;
            16'd7638: data <= 8'h00;
            16'd7639: data <= 8'hF8;
            16'd7640: data <= 8'hFF;
            16'd7641: data <= 8'hFF;
            16'd7642: data <= 8'h00;
            16'd7643: data <= 8'hF8;
            16'd7644: data <= 8'h00;
            16'd7645: data <= 8'hF8;
            16'd7646: data <= 8'h00;
            16'd7647: data <= 8'hF8;
            16'd7648: data <= 8'h00;
            16'd7649: data <= 8'hF8;
            16'd7650: data <= 8'h00;
            16'd7651: data <= 8'hF8;
            16'd7652: data <= 8'h00;
            16'd7653: data <= 8'hF8;
            16'd7654: data <= 8'h00;
            16'd7655: data <= 8'hF8;
            16'd7656: data <= 8'h00;
            16'd7657: data <= 8'hF8;
            16'd7658: data <= 8'h00;
            16'd7659: data <= 8'hF8;
            16'd7660: data <= 8'h00;
            16'd7661: data <= 8'hF8;
            16'd7662: data <= 8'h00;
            16'd7663: data <= 8'hF8;
            16'd7664: data <= 8'h00;
            16'd7665: data <= 8'hF8;
            16'd7666: data <= 8'h00;
            16'd7667: data <= 8'hF8;
            16'd7668: data <= 8'h00;
            16'd7669: data <= 8'hF8;
            16'd7670: data <= 8'h00;
            16'd7671: data <= 8'hF8;
            16'd7672: data <= 8'h00;
            16'd7673: data <= 8'hF8;
            16'd7674: data <= 8'h00;
            16'd7675: data <= 8'hF8;
            16'd7676: data <= 8'h00;
            16'd7677: data <= 8'hF8;
            16'd7678: data <= 8'h00;
            16'd7679: data <= 8'hF8;
            16'd7680: data <= 8'hFF;
            16'd7681: data <= 8'hFF;
            16'd7682: data <= 8'h00;
            16'd7683: data <= 8'hF8;
            16'd7684: data <= 8'h00;
            16'd7685: data <= 8'hF8;
            16'd7686: data <= 8'h00;
            16'd7687: data <= 8'hF8;
            16'd7688: data <= 8'h00;
            16'd7689: data <= 8'hF8;
            16'd7690: data <= 8'h00;
            16'd7691: data <= 8'hF8;
            16'd7692: data <= 8'h00;
            16'd7693: data <= 8'hF8;
            16'd7694: data <= 8'h00;
            16'd7695: data <= 8'hF8;
            16'd7696: data <= 8'h00;
            16'd7697: data <= 8'hF8;
            16'd7698: data <= 8'h00;
            16'd7699: data <= 8'hF8;
            16'd7700: data <= 8'h00;
            16'd7701: data <= 8'hF8;
            16'd7702: data <= 8'h00;
            16'd7703: data <= 8'hF8;
            16'd7704: data <= 8'h00;
            16'd7705: data <= 8'hF8;
            16'd7706: data <= 8'h00;
            16'd7707: data <= 8'hF8;
            16'd7708: data <= 8'h00;
            16'd7709: data <= 8'hF8;
            16'd7710: data <= 8'h00;
            16'd7711: data <= 8'hF8;
            16'd7712: data <= 8'h00;
            16'd7713: data <= 8'hF8;
            16'd7714: data <= 8'h00;
            16'd7715: data <= 8'hF8;
            16'd7716: data <= 8'h00;
            16'd7717: data <= 8'hF8;
            16'd7718: data <= 8'h00;
            16'd7719: data <= 8'hF8;
            16'd7720: data <= 8'hFF;
            16'd7721: data <= 8'hFF;
            16'd7722: data <= 8'h00;
            16'd7723: data <= 8'hF8;
            16'd7724: data <= 8'h00;
            16'd7725: data <= 8'hF8;
            16'd7726: data <= 8'h00;
            16'd7727: data <= 8'hF8;
            16'd7728: data <= 8'h00;
            16'd7729: data <= 8'hF8;
            16'd7730: data <= 8'h00;
            16'd7731: data <= 8'hF8;
            16'd7732: data <= 8'h00;
            16'd7733: data <= 8'hF8;
            16'd7734: data <= 8'h00;
            16'd7735: data <= 8'hF8;
            16'd7736: data <= 8'h00;
            16'd7737: data <= 8'hF8;
            16'd7738: data <= 8'h00;
            16'd7739: data <= 8'hF8;
            16'd7740: data <= 8'h00;
            16'd7741: data <= 8'hF8;
            16'd7742: data <= 8'h00;
            16'd7743: data <= 8'hF8;
            16'd7744: data <= 8'h00;
            16'd7745: data <= 8'hF8;
            16'd7746: data <= 8'h00;
            16'd7747: data <= 8'hF8;
            16'd7748: data <= 8'h00;
            16'd7749: data <= 8'hF8;
            16'd7750: data <= 8'h00;
            16'd7751: data <= 8'hF8;
            16'd7752: data <= 8'h00;
            16'd7753: data <= 8'hF8;
            16'd7754: data <= 8'h00;
            16'd7755: data <= 8'hF8;
            16'd7756: data <= 8'h00;
            16'd7757: data <= 8'hF8;
            16'd7758: data <= 8'h00;
            16'd7759: data <= 8'hF8;
            16'd7760: data <= 8'hFF;
            16'd7761: data <= 8'hFF;
            16'd7762: data <= 8'h00;
            16'd7763: data <= 8'hF8;
            16'd7764: data <= 8'h00;
            16'd7765: data <= 8'hF8;
            16'd7766: data <= 8'h00;
            16'd7767: data <= 8'hF8;
            16'd7768: data <= 8'h00;
            16'd7769: data <= 8'hF8;
            16'd7770: data <= 8'h00;
            16'd7771: data <= 8'hF8;
            16'd7772: data <= 8'h00;
            16'd7773: data <= 8'hF8;
            16'd7774: data <= 8'h00;
            16'd7775: data <= 8'hF8;
            16'd7776: data <= 8'h00;
            16'd7777: data <= 8'hF8;
            16'd7778: data <= 8'h00;
            16'd7779: data <= 8'hF8;
            16'd7780: data <= 8'h00;
            16'd7781: data <= 8'hF8;
            16'd7782: data <= 8'h00;
            16'd7783: data <= 8'hF8;
            16'd7784: data <= 8'h00;
            16'd7785: data <= 8'hF8;
            16'd7786: data <= 8'h00;
            16'd7787: data <= 8'hF8;
            16'd7788: data <= 8'h00;
            16'd7789: data <= 8'hF8;
            16'd7790: data <= 8'h00;
            16'd7791: data <= 8'hF8;
            16'd7792: data <= 8'h00;
            16'd7793: data <= 8'hF8;
            16'd7794: data <= 8'h00;
            16'd7795: data <= 8'hF8;
            16'd7796: data <= 8'h00;
            16'd7797: data <= 8'hF8;
            16'd7798: data <= 8'h00;
            16'd7799: data <= 8'hF8;
            16'd7800: data <= 8'hFF;
            16'd7801: data <= 8'hFF;
            16'd7802: data <= 8'h00;
            16'd7803: data <= 8'hF8;
            16'd7804: data <= 8'h00;
            16'd7805: data <= 8'hF8;
            16'd7806: data <= 8'h00;
            16'd7807: data <= 8'hF8;
            16'd7808: data <= 8'h00;
            16'd7809: data <= 8'hF8;
            16'd7810: data <= 8'h00;
            16'd7811: data <= 8'hF8;
            16'd7812: data <= 8'h00;
            16'd7813: data <= 8'hF8;
            16'd7814: data <= 8'h00;
            16'd7815: data <= 8'hF8;
            16'd7816: data <= 8'h00;
            16'd7817: data <= 8'hF8;
            16'd7818: data <= 8'h00;
            16'd7819: data <= 8'hF8;
            16'd7820: data <= 8'h00;
            16'd7821: data <= 8'hF8;
            16'd7822: data <= 8'h00;
            16'd7823: data <= 8'hF8;
            16'd7824: data <= 8'h00;
            16'd7825: data <= 8'hF8;
            16'd7826: data <= 8'h00;
            16'd7827: data <= 8'hF8;
            16'd7828: data <= 8'h00;
            16'd7829: data <= 8'hF8;
            16'd7830: data <= 8'h00;
            16'd7831: data <= 8'hF8;
            16'd7832: data <= 8'h00;
            16'd7833: data <= 8'hF8;
            16'd7834: data <= 8'h00;
            16'd7835: data <= 8'hF8;
            16'd7836: data <= 8'h00;
            16'd7837: data <= 8'hF8;
            16'd7838: data <= 8'h00;
            16'd7839: data <= 8'hF8;
            16'd7840: data <= 8'hFF;
            16'd7841: data <= 8'hFF;
            16'd7842: data <= 8'h00;
            16'd7843: data <= 8'hF8;
            16'd7844: data <= 8'h00;
            16'd7845: data <= 8'hF8;
            16'd7846: data <= 8'h00;
            16'd7847: data <= 8'hF8;
            16'd7848: data <= 8'h00;
            16'd7849: data <= 8'hF8;
            16'd7850: data <= 8'h00;
            16'd7851: data <= 8'hF8;
            16'd7852: data <= 8'h00;
            16'd7853: data <= 8'hF8;
            16'd7854: data <= 8'h00;
            16'd7855: data <= 8'hF8;
            16'd7856: data <= 8'h00;
            16'd7857: data <= 8'hF8;
            16'd7858: data <= 8'h00;
            16'd7859: data <= 8'hF8;
            16'd7860: data <= 8'h00;
            16'd7861: data <= 8'hF8;
            16'd7862: data <= 8'h00;
            16'd7863: data <= 8'hF8;
            16'd7864: data <= 8'h00;
            16'd7865: data <= 8'hF8;
            16'd7866: data <= 8'h00;
            16'd7867: data <= 8'hF8;
            16'd7868: data <= 8'h00;
            16'd7869: data <= 8'hF8;
            16'd7870: data <= 8'h00;
            16'd7871: data <= 8'hF8;
            16'd7872: data <= 8'h00;
            16'd7873: data <= 8'hF8;
            16'd7874: data <= 8'h00;
            16'd7875: data <= 8'hF8;
            16'd7876: data <= 8'h00;
            16'd7877: data <= 8'hF8;
            16'd7878: data <= 8'h00;
            16'd7879: data <= 8'hF8;
            16'd7880: data <= 8'hFF;
            16'd7881: data <= 8'hFF;
            16'd7882: data <= 8'h00;
            16'd7883: data <= 8'hF8;
            16'd7884: data <= 8'h00;
            16'd7885: data <= 8'hF8;
            16'd7886: data <= 8'h00;
            16'd7887: data <= 8'hF8;
            16'd7888: data <= 8'h00;
            16'd7889: data <= 8'hF8;
            16'd7890: data <= 8'h00;
            16'd7891: data <= 8'hF8;
            16'd7892: data <= 8'h00;
            16'd7893: data <= 8'hF8;
            16'd7894: data <= 8'h00;
            16'd7895: data <= 8'hF8;
            16'd7896: data <= 8'h00;
            16'd7897: data <= 8'hF8;
            16'd7898: data <= 8'h00;
            16'd7899: data <= 8'hF8;
            16'd7900: data <= 8'h00;
            16'd7901: data <= 8'hF8;
            16'd7902: data <= 8'h00;
            16'd7903: data <= 8'hF8;
            16'd7904: data <= 8'h00;
            16'd7905: data <= 8'hF8;
            16'd7906: data <= 8'h00;
            16'd7907: data <= 8'hF8;
            16'd7908: data <= 8'h00;
            16'd7909: data <= 8'hF8;
            16'd7910: data <= 8'h00;
            16'd7911: data <= 8'hF8;
            16'd7912: data <= 8'h00;
            16'd7913: data <= 8'hF8;
            16'd7914: data <= 8'h00;
            16'd7915: data <= 8'hF8;
            16'd7916: data <= 8'h00;
            16'd7917: data <= 8'hF8;
            16'd7918: data <= 8'h00;
            16'd7919: data <= 8'hF8;
            16'd7920: data <= 8'hFF;
            16'd7921: data <= 8'hFF;
            16'd7922: data <= 8'h00;
            16'd7923: data <= 8'hF8;
            16'd7924: data <= 8'h00;
            16'd7925: data <= 8'hF8;
            16'd7926: data <= 8'h00;
            16'd7927: data <= 8'hF8;
            16'd7928: data <= 8'h00;
            16'd7929: data <= 8'hF8;
            16'd7930: data <= 8'h00;
            16'd7931: data <= 8'hF8;
            16'd7932: data <= 8'h00;
            16'd7933: data <= 8'hF8;
            16'd7934: data <= 8'h00;
            16'd7935: data <= 8'hF8;
            16'd7936: data <= 8'h00;
            16'd7937: data <= 8'hF8;
            16'd7938: data <= 8'h00;
            16'd7939: data <= 8'hF8;
            16'd7940: data <= 8'h00;
            16'd7941: data <= 8'hF8;
            16'd7942: data <= 8'h00;
            16'd7943: data <= 8'hF8;
            16'd7944: data <= 8'h00;
            16'd7945: data <= 8'hF8;
            16'd7946: data <= 8'h00;
            16'd7947: data <= 8'hF8;
            16'd7948: data <= 8'h00;
            16'd7949: data <= 8'hF8;
            16'd7950: data <= 8'h00;
            16'd7951: data <= 8'hF8;
            16'd7952: data <= 8'h00;
            16'd7953: data <= 8'hF8;
            16'd7954: data <= 8'h00;
            16'd7955: data <= 8'hF8;
            16'd7956: data <= 8'h00;
            16'd7957: data <= 8'hF8;
            16'd7958: data <= 8'h00;
            16'd7959: data <= 8'hF8;
            16'd7960: data <= 8'hFF;
            16'd7961: data <= 8'hFF;
            16'd7962: data <= 8'h00;
            16'd7963: data <= 8'hF8;
            16'd7964: data <= 8'h00;
            16'd7965: data <= 8'hF8;
            16'd7966: data <= 8'h00;
            16'd7967: data <= 8'hF8;
            16'd7968: data <= 8'h00;
            16'd7969: data <= 8'hF8;
            16'd7970: data <= 8'h00;
            16'd7971: data <= 8'hF8;
            16'd7972: data <= 8'h00;
            16'd7973: data <= 8'hF8;
            16'd7974: data <= 8'h00;
            16'd7975: data <= 8'hF8;
            16'd7976: data <= 8'h00;
            16'd7977: data <= 8'hF8;
            16'd7978: data <= 8'h00;
            16'd7979: data <= 8'hF8;
            16'd7980: data <= 8'h00;
            16'd7981: data <= 8'hF8;
            16'd7982: data <= 8'h00;
            16'd7983: data <= 8'hF8;
            16'd7984: data <= 8'h00;
            16'd7985: data <= 8'hF8;
            16'd7986: data <= 8'h00;
            16'd7987: data <= 8'hF8;
            16'd7988: data <= 8'h00;
            16'd7989: data <= 8'hF8;
            16'd7990: data <= 8'h00;
            16'd7991: data <= 8'hF8;
            16'd7992: data <= 8'h00;
            16'd7993: data <= 8'hF8;
            16'd7994: data <= 8'h00;
            16'd7995: data <= 8'hF8;
            16'd7996: data <= 8'h00;
            16'd7997: data <= 8'hF8;
            16'd7998: data <= 8'h00;
            16'd7999: data <= 8'hF8;
            16'd8000: data <= 8'hFF;
            16'd8001: data <= 8'hFF;
            16'd8002: data <= 8'h00;
            16'd8003: data <= 8'hF8;
            16'd8004: data <= 8'h00;
            16'd8005: data <= 8'hF8;
            16'd8006: data <= 8'h00;
            16'd8007: data <= 8'hF8;
            16'd8008: data <= 8'h00;
            16'd8009: data <= 8'hF8;
            16'd8010: data <= 8'h00;
            16'd8011: data <= 8'hF8;
            16'd8012: data <= 8'h00;
            16'd8013: data <= 8'hF8;
            16'd8014: data <= 8'h00;
            16'd8015: data <= 8'hF8;
            16'd8016: data <= 8'h00;
            16'd8017: data <= 8'hF8;
            16'd8018: data <= 8'h00;
            16'd8019: data <= 8'hF8;
            16'd8020: data <= 8'h00;
            16'd8021: data <= 8'hF8;
            16'd8022: data <= 8'h00;
            16'd8023: data <= 8'hF8;
            16'd8024: data <= 8'h00;
            16'd8025: data <= 8'hF8;
            16'd8026: data <= 8'h00;
            16'd8027: data <= 8'hF8;
            16'd8028: data <= 8'h00;
            16'd8029: data <= 8'hF8;
            16'd8030: data <= 8'h00;
            16'd8031: data <= 8'hF8;
            16'd8032: data <= 8'h00;
            16'd8033: data <= 8'hF8;
            16'd8034: data <= 8'h00;
            16'd8035: data <= 8'hF8;
            16'd8036: data <= 8'h00;
            16'd8037: data <= 8'hF8;
            16'd8038: data <= 8'h00;
            16'd8039: data <= 8'hF8;
            16'd8040: data <= 8'hFF;
            16'd8041: data <= 8'hFF;
            16'd8042: data <= 8'h00;
            16'd8043: data <= 8'hF8;
            16'd8044: data <= 8'h00;
            16'd8045: data <= 8'hF8;
            16'd8046: data <= 8'h00;
            16'd8047: data <= 8'hF8;
            16'd8048: data <= 8'h00;
            16'd8049: data <= 8'hF8;
            16'd8050: data <= 8'h00;
            16'd8051: data <= 8'hF8;
            16'd8052: data <= 8'h00;
            16'd8053: data <= 8'hF8;
            16'd8054: data <= 8'h00;
            16'd8055: data <= 8'hF8;
            16'd8056: data <= 8'h00;
            16'd8057: data <= 8'hF8;
            16'd8058: data <= 8'h00;
            16'd8059: data <= 8'hF8;
            16'd8060: data <= 8'h00;
            16'd8061: data <= 8'hF8;
            16'd8062: data <= 8'h00;
            16'd8063: data <= 8'hF8;
            16'd8064: data <= 8'h00;
            16'd8065: data <= 8'hF8;
            16'd8066: data <= 8'h00;
            16'd8067: data <= 8'hF8;
            16'd8068: data <= 8'h00;
            16'd8069: data <= 8'hF8;
            16'd8070: data <= 8'h00;
            16'd8071: data <= 8'hF8;
            16'd8072: data <= 8'h00;
            16'd8073: data <= 8'hF8;
            16'd8074: data <= 8'h00;
            16'd8075: data <= 8'hF8;
            16'd8076: data <= 8'h00;
            16'd8077: data <= 8'hF8;
            16'd8078: data <= 8'h00;
            16'd8079: data <= 8'hF8;
            16'd8080: data <= 8'hFF;
            16'd8081: data <= 8'hFF;
            16'd8082: data <= 8'h00;
            16'd8083: data <= 8'hF8;
            16'd8084: data <= 8'h00;
            16'd8085: data <= 8'hF8;
            16'd8086: data <= 8'h00;
            16'd8087: data <= 8'hF8;
            16'd8088: data <= 8'h00;
            16'd8089: data <= 8'hF8;
            16'd8090: data <= 8'h00;
            16'd8091: data <= 8'hF8;
            16'd8092: data <= 8'h00;
            16'd8093: data <= 8'hF8;
            16'd8094: data <= 8'h00;
            16'd8095: data <= 8'hF8;
            16'd8096: data <= 8'h00;
            16'd8097: data <= 8'hF8;
            16'd8098: data <= 8'h00;
            16'd8099: data <= 8'hF8;
            16'd8100: data <= 8'h00;
            16'd8101: data <= 8'hF8;
            16'd8102: data <= 8'h00;
            16'd8103: data <= 8'hF8;
            16'd8104: data <= 8'h00;
            16'd8105: data <= 8'hF8;
            16'd8106: data <= 8'h00;
            16'd8107: data <= 8'hF8;
            16'd8108: data <= 8'h00;
            16'd8109: data <= 8'hF8;
            16'd8110: data <= 8'h00;
            16'd8111: data <= 8'hF8;
            16'd8112: data <= 8'h00;
            16'd8113: data <= 8'hF8;
            16'd8114: data <= 8'h00;
            16'd8115: data <= 8'hF8;
            16'd8116: data <= 8'h00;
            16'd8117: data <= 8'hF8;
            16'd8118: data <= 8'h00;
            16'd8119: data <= 8'hF8;
            16'd8120: data <= 8'hFF;
            16'd8121: data <= 8'hFF;
            16'd8122: data <= 8'h00;
            16'd8123: data <= 8'hF8;
            16'd8124: data <= 8'h00;
            16'd8125: data <= 8'hF8;
            16'd8126: data <= 8'h00;
            16'd8127: data <= 8'hF8;
            16'd8128: data <= 8'h00;
            16'd8129: data <= 8'hF8;
            16'd8130: data <= 8'h00;
            16'd8131: data <= 8'hF8;
            16'd8132: data <= 8'h00;
            16'd8133: data <= 8'hF8;
            16'd8134: data <= 8'h00;
            16'd8135: data <= 8'hF8;
            16'd8136: data <= 8'h00;
            16'd8137: data <= 8'hF8;
            16'd8138: data <= 8'h00;
            16'd8139: data <= 8'hF8;
            16'd8140: data <= 8'h00;
            16'd8141: data <= 8'hF8;
            16'd8142: data <= 8'h00;
            16'd8143: data <= 8'hF8;
            16'd8144: data <= 8'h00;
            16'd8145: data <= 8'hF8;
            16'd8146: data <= 8'h00;
            16'd8147: data <= 8'hF8;
            16'd8148: data <= 8'h00;
            16'd8149: data <= 8'hF8;
            16'd8150: data <= 8'h00;
            16'd8151: data <= 8'hF8;
            16'd8152: data <= 8'h00;
            16'd8153: data <= 8'hF8;
            16'd8154: data <= 8'h00;
            16'd8155: data <= 8'hF8;
            16'd8156: data <= 8'h00;
            16'd8157: data <= 8'hF8;
            16'd8158: data <= 8'h00;
            16'd8159: data <= 8'hF8;
            16'd8160: data <= 8'hFF;
            16'd8161: data <= 8'hFF;
            16'd8162: data <= 8'h00;
            16'd8163: data <= 8'hF8;
            16'd8164: data <= 8'h00;
            16'd8165: data <= 8'hF8;
            16'd8166: data <= 8'h00;
            16'd8167: data <= 8'hF8;
            16'd8168: data <= 8'h00;
            16'd8169: data <= 8'hF8;
            16'd8170: data <= 8'h00;
            16'd8171: data <= 8'hF8;
            16'd8172: data <= 8'h00;
            16'd8173: data <= 8'hF8;
            16'd8174: data <= 8'h00;
            16'd8175: data <= 8'hF8;
            16'd8176: data <= 8'h00;
            16'd8177: data <= 8'hF8;
            16'd8178: data <= 8'h00;
            16'd8179: data <= 8'hF8;
            16'd8180: data <= 8'h00;
            16'd8181: data <= 8'hF8;
            16'd8182: data <= 8'h00;
            16'd8183: data <= 8'hF8;
            16'd8184: data <= 8'h00;
            16'd8185: data <= 8'hF8;
            16'd8186: data <= 8'h00;
            16'd8187: data <= 8'hF8;
            16'd8188: data <= 8'h00;
            16'd8189: data <= 8'hF8;
            16'd8190: data <= 8'h00;
            16'd8191: data <= 8'hF8;
            16'd8192: data <= 8'h00;
            16'd8193: data <= 8'hF8;
            16'd8194: data <= 8'h00;
            16'd8195: data <= 8'hF8;
            16'd8196: data <= 8'h00;
            16'd8197: data <= 8'hF8;
            16'd8198: data <= 8'h00;
            16'd8199: data <= 8'hF8;
            16'd8200: data <= 8'hFF;
            16'd8201: data <= 8'hFF;
            16'd8202: data <= 8'h00;
            16'd8203: data <= 8'hF8;
            16'd8204: data <= 8'h00;
            16'd8205: data <= 8'hF8;
            16'd8206: data <= 8'h00;
            16'd8207: data <= 8'hF8;
            16'd8208: data <= 8'h00;
            16'd8209: data <= 8'hF8;
            16'd8210: data <= 8'h00;
            16'd8211: data <= 8'hF8;
            16'd8212: data <= 8'h00;
            16'd8213: data <= 8'hF8;
            16'd8214: data <= 8'h00;
            16'd8215: data <= 8'hF8;
            16'd8216: data <= 8'h00;
            16'd8217: data <= 8'hF8;
            16'd8218: data <= 8'h00;
            16'd8219: data <= 8'hF8;
            16'd8220: data <= 8'h00;
            16'd8221: data <= 8'hF8;
            16'd8222: data <= 8'h00;
            16'd8223: data <= 8'hF8;
            16'd8224: data <= 8'h00;
            16'd8225: data <= 8'hF8;
            16'd8226: data <= 8'h00;
            16'd8227: data <= 8'hF8;
            16'd8228: data <= 8'h00;
            16'd8229: data <= 8'hF8;
            16'd8230: data <= 8'h00;
            16'd8231: data <= 8'hF8;
            16'd8232: data <= 8'h00;
            16'd8233: data <= 8'hF8;
            16'd8234: data <= 8'h00;
            16'd8235: data <= 8'hF8;
            16'd8236: data <= 8'h00;
            16'd8237: data <= 8'hF8;
            16'd8238: data <= 8'h00;
            16'd8239: data <= 8'hF8;
            16'd8240: data <= 8'hFF;
            16'd8241: data <= 8'hFF;
            16'd8242: data <= 8'h00;
            16'd8243: data <= 8'hF8;
            16'd8244: data <= 8'h00;
            16'd8245: data <= 8'hF8;
            16'd8246: data <= 8'h00;
            16'd8247: data <= 8'hF8;
            16'd8248: data <= 8'h00;
            16'd8249: data <= 8'hF8;
            16'd8250: data <= 8'h00;
            16'd8251: data <= 8'hF8;
            16'd8252: data <= 8'h00;
            16'd8253: data <= 8'hF8;
            16'd8254: data <= 8'h00;
            16'd8255: data <= 8'hF8;
            16'd8256: data <= 8'h00;
            16'd8257: data <= 8'hF8;
            16'd8258: data <= 8'h00;
            16'd8259: data <= 8'hF8;
            16'd8260: data <= 8'h00;
            16'd8261: data <= 8'hF8;
            16'd8262: data <= 8'h00;
            16'd8263: data <= 8'hF8;
            16'd8264: data <= 8'h00;
            16'd8265: data <= 8'hF8;
            16'd8266: data <= 8'h00;
            16'd8267: data <= 8'hF8;
            16'd8268: data <= 8'h00;
            16'd8269: data <= 8'hF8;
            16'd8270: data <= 8'h00;
            16'd8271: data <= 8'hF8;
            16'd8272: data <= 8'h00;
            16'd8273: data <= 8'hF8;
            16'd8274: data <= 8'h00;
            16'd8275: data <= 8'hF8;
            16'd8276: data <= 8'h00;
            16'd8277: data <= 8'hF8;
            16'd8278: data <= 8'h00;
            16'd8279: data <= 8'hF8;
            16'd8280: data <= 8'hFF;
            16'd8281: data <= 8'hFF;
            16'd8282: data <= 8'h00;
            16'd8283: data <= 8'hF8;
            16'd8284: data <= 8'h00;
            16'd8285: data <= 8'hF8;
            16'd8286: data <= 8'h00;
            16'd8287: data <= 8'hF8;
            16'd8288: data <= 8'h00;
            16'd8289: data <= 8'hF8;
            16'd8290: data <= 8'h00;
            16'd8291: data <= 8'hF8;
            16'd8292: data <= 8'h00;
            16'd8293: data <= 8'hF8;
            16'd8294: data <= 8'h00;
            16'd8295: data <= 8'hF8;
            16'd8296: data <= 8'h00;
            16'd8297: data <= 8'hF8;
            16'd8298: data <= 8'h00;
            16'd8299: data <= 8'hF8;
            16'd8300: data <= 8'h00;
            16'd8301: data <= 8'hF8;
            16'd8302: data <= 8'h00;
            16'd8303: data <= 8'hF8;
            16'd8304: data <= 8'h00;
            16'd8305: data <= 8'hF8;
            16'd8306: data <= 8'h00;
            16'd8307: data <= 8'hF8;
            16'd8308: data <= 8'h00;
            16'd8309: data <= 8'hF8;
            16'd8310: data <= 8'h00;
            16'd8311: data <= 8'hF8;
            16'd8312: data <= 8'h00;
            16'd8313: data <= 8'hF8;
            16'd8314: data <= 8'h00;
            16'd8315: data <= 8'hF8;
            16'd8316: data <= 8'h00;
            16'd8317: data <= 8'hF8;
            16'd8318: data <= 8'h00;
            16'd8319: data <= 8'hF8;
            16'd8320: data <= 8'hFF;
            16'd8321: data <= 8'hFF;
            16'd8322: data <= 8'h00;
            16'd8323: data <= 8'hF8;
            16'd8324: data <= 8'h00;
            16'd8325: data <= 8'hF8;
            16'd8326: data <= 8'h00;
            16'd8327: data <= 8'hF8;
            16'd8328: data <= 8'h00;
            16'd8329: data <= 8'hF8;
            16'd8330: data <= 8'h00;
            16'd8331: data <= 8'hF8;
            16'd8332: data <= 8'h00;
            16'd8333: data <= 8'hF8;
            16'd8334: data <= 8'h00;
            16'd8335: data <= 8'hF8;
            16'd8336: data <= 8'h00;
            16'd8337: data <= 8'hF8;
            16'd8338: data <= 8'h00;
            16'd8339: data <= 8'hF8;
            16'd8340: data <= 8'h00;
            16'd8341: data <= 8'hF8;
            16'd8342: data <= 8'h00;
            16'd8343: data <= 8'hF8;
            16'd8344: data <= 8'h00;
            16'd8345: data <= 8'hF8;
            16'd8346: data <= 8'h00;
            16'd8347: data <= 8'hF8;
            16'd8348: data <= 8'h00;
            16'd8349: data <= 8'hF8;
            16'd8350: data <= 8'h00;
            16'd8351: data <= 8'hF8;
            16'd8352: data <= 8'h00;
            16'd8353: data <= 8'hF8;
            16'd8354: data <= 8'h00;
            16'd8355: data <= 8'hF8;
            16'd8356: data <= 8'h00;
            16'd8357: data <= 8'hF8;
            16'd8358: data <= 8'h00;
            16'd8359: data <= 8'hF8;
            16'd8360: data <= 8'hFF;
            16'd8361: data <= 8'hFF;
            16'd8362: data <= 8'h00;
            16'd8363: data <= 8'hF8;
            16'd8364: data <= 8'h00;
            16'd8365: data <= 8'hF8;
            16'd8366: data <= 8'h00;
            16'd8367: data <= 8'hF8;
            16'd8368: data <= 8'h00;
            16'd8369: data <= 8'hF8;
            16'd8370: data <= 8'h00;
            16'd8371: data <= 8'hF8;
            16'd8372: data <= 8'h00;
            16'd8373: data <= 8'hF8;
            16'd8374: data <= 8'h00;
            16'd8375: data <= 8'hF8;
            16'd8376: data <= 8'h00;
            16'd8377: data <= 8'hF8;
            16'd8378: data <= 8'h00;
            16'd8379: data <= 8'hF8;
            16'd8380: data <= 8'h00;
            16'd8381: data <= 8'hF8;
            16'd8382: data <= 8'h00;
            16'd8383: data <= 8'hF8;
            16'd8384: data <= 8'h00;
            16'd8385: data <= 8'hF8;
            16'd8386: data <= 8'h00;
            16'd8387: data <= 8'hF8;
            16'd8388: data <= 8'h00;
            16'd8389: data <= 8'hF8;
            16'd8390: data <= 8'h00;
            16'd8391: data <= 8'hF8;
            16'd8392: data <= 8'h00;
            16'd8393: data <= 8'hF8;
            16'd8394: data <= 8'h00;
            16'd8395: data <= 8'hF8;
            16'd8396: data <= 8'h00;
            16'd8397: data <= 8'hF8;
            16'd8398: data <= 8'h00;
            16'd8399: data <= 8'hF8;
            16'd8400: data <= 8'hFF;
            16'd8401: data <= 8'hFF;
            16'd8402: data <= 8'h00;
            16'd8403: data <= 8'hF8;
            16'd8404: data <= 8'h00;
            16'd8405: data <= 8'hF8;
            16'd8406: data <= 8'h00;
            16'd8407: data <= 8'hF8;
            16'd8408: data <= 8'h00;
            16'd8409: data <= 8'hF8;
            16'd8410: data <= 8'h00;
            16'd8411: data <= 8'hF8;
            16'd8412: data <= 8'h00;
            16'd8413: data <= 8'hF8;
            16'd8414: data <= 8'h00;
            16'd8415: data <= 8'hF8;
            16'd8416: data <= 8'h00;
            16'd8417: data <= 8'hF8;
            16'd8418: data <= 8'h00;
            16'd8419: data <= 8'hF8;
            16'd8420: data <= 8'h00;
            16'd8421: data <= 8'hF8;
            16'd8422: data <= 8'h00;
            16'd8423: data <= 8'hF8;
            16'd8424: data <= 8'h00;
            16'd8425: data <= 8'hF8;
            16'd8426: data <= 8'h00;
            16'd8427: data <= 8'hF8;
            16'd8428: data <= 8'h00;
            16'd8429: data <= 8'hF8;
            16'd8430: data <= 8'h00;
            16'd8431: data <= 8'hF8;
            16'd8432: data <= 8'h00;
            16'd8433: data <= 8'hF8;
            16'd8434: data <= 8'h00;
            16'd8435: data <= 8'hF8;
            16'd8436: data <= 8'h00;
            16'd8437: data <= 8'hF8;
            16'd8438: data <= 8'h00;
            16'd8439: data <= 8'hF8;
            16'd8440: data <= 8'hFF;
            16'd8441: data <= 8'hFF;
            16'd8442: data <= 8'h00;
            16'd8443: data <= 8'hF8;
            16'd8444: data <= 8'h00;
            16'd8445: data <= 8'hF8;
            16'd8446: data <= 8'h00;
            16'd8447: data <= 8'hF8;
            16'd8448: data <= 8'h00;
            16'd8449: data <= 8'hF8;
            16'd8450: data <= 8'h00;
            16'd8451: data <= 8'hF8;
            16'd8452: data <= 8'h00;
            16'd8453: data <= 8'hF8;
            16'd8454: data <= 8'h00;
            16'd8455: data <= 8'hF8;
            16'd8456: data <= 8'h00;
            16'd8457: data <= 8'hF8;
            16'd8458: data <= 8'h00;
            16'd8459: data <= 8'hF8;
            16'd8460: data <= 8'h00;
            16'd8461: data <= 8'hF8;
            16'd8462: data <= 8'h00;
            16'd8463: data <= 8'hF8;
            16'd8464: data <= 8'h00;
            16'd8465: data <= 8'hF8;
            16'd8466: data <= 8'h00;
            16'd8467: data <= 8'hF8;
            16'd8468: data <= 8'h00;
            16'd8469: data <= 8'hF8;
            16'd8470: data <= 8'h00;
            16'd8471: data <= 8'hF8;
            16'd8472: data <= 8'h00;
            16'd8473: data <= 8'hF8;
            16'd8474: data <= 8'h00;
            16'd8475: data <= 8'hF8;
            16'd8476: data <= 8'h00;
            16'd8477: data <= 8'hF8;
            16'd8478: data <= 8'h00;
            16'd8479: data <= 8'hF8;
            16'd8480: data <= 8'hFF;
            16'd8481: data <= 8'hFF;
            16'd8482: data <= 8'h00;
            16'd8483: data <= 8'hF8;
            16'd8484: data <= 8'h00;
            16'd8485: data <= 8'hF8;
            16'd8486: data <= 8'h00;
            16'd8487: data <= 8'hF8;
            16'd8488: data <= 8'h00;
            16'd8489: data <= 8'hF8;
            16'd8490: data <= 8'h00;
            16'd8491: data <= 8'hF8;
            16'd8492: data <= 8'h00;
            16'd8493: data <= 8'hF8;
            16'd8494: data <= 8'h00;
            16'd8495: data <= 8'hF8;
            16'd8496: data <= 8'h00;
            16'd8497: data <= 8'hF8;
            16'd8498: data <= 8'h00;
            16'd8499: data <= 8'hF8;
            16'd8500: data <= 8'h00;
            16'd8501: data <= 8'hF8;
            16'd8502: data <= 8'h00;
            16'd8503: data <= 8'hF8;
            16'd8504: data <= 8'h00;
            16'd8505: data <= 8'hF8;
            16'd8506: data <= 8'h00;
            16'd8507: data <= 8'hF8;
            16'd8508: data <= 8'h00;
            16'd8509: data <= 8'hF8;
            16'd8510: data <= 8'h00;
            16'd8511: data <= 8'hF8;
            16'd8512: data <= 8'h00;
            16'd8513: data <= 8'hF8;
            16'd8514: data <= 8'h00;
            16'd8515: data <= 8'hF8;
            16'd8516: data <= 8'h00;
            16'd8517: data <= 8'hF8;
            16'd8518: data <= 8'h00;
            16'd8519: data <= 8'hF8;
            16'd8520: data <= 8'hFF;
            16'd8521: data <= 8'hFF;
            16'd8522: data <= 8'h00;
            16'd8523: data <= 8'hF8;
            16'd8524: data <= 8'h00;
            16'd8525: data <= 8'hF8;
            16'd8526: data <= 8'h00;
            16'd8527: data <= 8'hF8;
            16'd8528: data <= 8'h00;
            16'd8529: data <= 8'hF8;
            16'd8530: data <= 8'h00;
            16'd8531: data <= 8'hF8;
            16'd8532: data <= 8'h00;
            16'd8533: data <= 8'hF8;
            16'd8534: data <= 8'h00;
            16'd8535: data <= 8'hF8;
            16'd8536: data <= 8'h00;
            16'd8537: data <= 8'hF8;
            16'd8538: data <= 8'h00;
            16'd8539: data <= 8'hF8;
            16'd8540: data <= 8'h00;
            16'd8541: data <= 8'hF8;
            16'd8542: data <= 8'h00;
            16'd8543: data <= 8'hF8;
            16'd8544: data <= 8'h00;
            16'd8545: data <= 8'hF8;
            16'd8546: data <= 8'h00;
            16'd8547: data <= 8'hF8;
            16'd8548: data <= 8'h00;
            16'd8549: data <= 8'hF8;
            16'd8550: data <= 8'h00;
            16'd8551: data <= 8'hF8;
            16'd8552: data <= 8'h00;
            16'd8553: data <= 8'hF8;
            16'd8554: data <= 8'h00;
            16'd8555: data <= 8'hF8;
            16'd8556: data <= 8'h00;
            16'd8557: data <= 8'hF8;
            16'd8558: data <= 8'h00;
            16'd8559: data <= 8'hF8;
            16'd8560: data <= 8'hFF;
            16'd8561: data <= 8'hFF;
            16'd8562: data <= 8'h00;
            16'd8563: data <= 8'hF8;
            16'd8564: data <= 8'h00;
            16'd8565: data <= 8'hF8;
            16'd8566: data <= 8'h00;
            16'd8567: data <= 8'hF8;
            16'd8568: data <= 8'h00;
            16'd8569: data <= 8'hF8;
            16'd8570: data <= 8'h00;
            16'd8571: data <= 8'hF8;
            16'd8572: data <= 8'h00;
            16'd8573: data <= 8'hF8;
            16'd8574: data <= 8'h00;
            16'd8575: data <= 8'hF8;
            16'd8576: data <= 8'h00;
            16'd8577: data <= 8'hF8;
            16'd8578: data <= 8'h00;
            16'd8579: data <= 8'hF8;
            16'd8580: data <= 8'h00;
            16'd8581: data <= 8'hF8;
            16'd8582: data <= 8'h00;
            16'd8583: data <= 8'hF8;
            16'd8584: data <= 8'h00;
            16'd8585: data <= 8'hF8;
            16'd8586: data <= 8'h00;
            16'd8587: data <= 8'hF8;
            16'd8588: data <= 8'h00;
            16'd8589: data <= 8'hF8;
            16'd8590: data <= 8'h00;
            16'd8591: data <= 8'hF8;
            16'd8592: data <= 8'h00;
            16'd8593: data <= 8'hF8;
            16'd8594: data <= 8'h00;
            16'd8595: data <= 8'hF8;
            16'd8596: data <= 8'h00;
            16'd8597: data <= 8'hF8;
            16'd8598: data <= 8'h00;
            16'd8599: data <= 8'hF8;
            16'd8600: data <= 8'hFF;
            16'd8601: data <= 8'hFF;
            16'd8602: data <= 8'h00;
            16'd8603: data <= 8'hF8;
            16'd8604: data <= 8'h00;
            16'd8605: data <= 8'hF8;
            16'd8606: data <= 8'h00;
            16'd8607: data <= 8'hF8;
            16'd8608: data <= 8'h00;
            16'd8609: data <= 8'hF8;
            16'd8610: data <= 8'h00;
            16'd8611: data <= 8'hF8;
            16'd8612: data <= 8'h00;
            16'd8613: data <= 8'hF8;
            16'd8614: data <= 8'h00;
            16'd8615: data <= 8'hF8;
            16'd8616: data <= 8'h00;
            16'd8617: data <= 8'hF8;
            16'd8618: data <= 8'h00;
            16'd8619: data <= 8'hF8;
            16'd8620: data <= 8'h00;
            16'd8621: data <= 8'hF8;
            16'd8622: data <= 8'h00;
            16'd8623: data <= 8'hF8;
            16'd8624: data <= 8'h00;
            16'd8625: data <= 8'hF8;
            16'd8626: data <= 8'h00;
            16'd8627: data <= 8'hF8;
            16'd8628: data <= 8'h00;
            16'd8629: data <= 8'hF8;
            16'd8630: data <= 8'h00;
            16'd8631: data <= 8'hF8;
            16'd8632: data <= 8'h00;
            16'd8633: data <= 8'hF8;
            16'd8634: data <= 8'h00;
            16'd8635: data <= 8'hF8;
            16'd8636: data <= 8'h00;
            16'd8637: data <= 8'hF8;
            16'd8638: data <= 8'h00;
            16'd8639: data <= 8'hF8;
            16'd8640: data <= 8'hFF;
            16'd8641: data <= 8'hFF;
            16'd8642: data <= 8'h00;
            16'd8643: data <= 8'hF8;
            16'd8644: data <= 8'h00;
            16'd8645: data <= 8'hF8;
            16'd8646: data <= 8'h00;
            16'd8647: data <= 8'hF8;
            16'd8648: data <= 8'h00;
            16'd8649: data <= 8'hF8;
            16'd8650: data <= 8'h00;
            16'd8651: data <= 8'hF8;
            16'd8652: data <= 8'h00;
            16'd8653: data <= 8'hF8;
            16'd8654: data <= 8'h00;
            16'd8655: data <= 8'hF8;
            16'd8656: data <= 8'h00;
            16'd8657: data <= 8'hF8;
            16'd8658: data <= 8'h00;
            16'd8659: data <= 8'hF8;
            16'd8660: data <= 8'h00;
            16'd8661: data <= 8'hF8;
            16'd8662: data <= 8'h00;
            16'd8663: data <= 8'hF8;
            16'd8664: data <= 8'h00;
            16'd8665: data <= 8'hF8;
            16'd8666: data <= 8'h00;
            16'd8667: data <= 8'hF8;
            16'd8668: data <= 8'h00;
            16'd8669: data <= 8'hF8;
            16'd8670: data <= 8'h00;
            16'd8671: data <= 8'hF8;
            16'd8672: data <= 8'h00;
            16'd8673: data <= 8'hF8;
            16'd8674: data <= 8'h00;
            16'd8675: data <= 8'hF8;
            16'd8676: data <= 8'h00;
            16'd8677: data <= 8'hF8;
            16'd8678: data <= 8'h00;
            16'd8679: data <= 8'hF8;
            16'd8680: data <= 8'hFF;
            16'd8681: data <= 8'hFF;
            16'd8682: data <= 8'h00;
            16'd8683: data <= 8'hF8;
            16'd8684: data <= 8'h00;
            16'd8685: data <= 8'hF8;
            16'd8686: data <= 8'h00;
            16'd8687: data <= 8'hF8;
            16'd8688: data <= 8'h00;
            16'd8689: data <= 8'hF8;
            16'd8690: data <= 8'h00;
            16'd8691: data <= 8'hF8;
            16'd8692: data <= 8'h00;
            16'd8693: data <= 8'hF8;
            16'd8694: data <= 8'h00;
            16'd8695: data <= 8'hF8;
            16'd8696: data <= 8'h00;
            16'd8697: data <= 8'hF8;
            16'd8698: data <= 8'h00;
            16'd8699: data <= 8'hF8;
            16'd8700: data <= 8'h00;
            16'd8701: data <= 8'hF8;
            16'd8702: data <= 8'h00;
            16'd8703: data <= 8'hF8;
            16'd8704: data <= 8'h00;
            16'd8705: data <= 8'hF8;
            16'd8706: data <= 8'h00;
            16'd8707: data <= 8'hF8;
            16'd8708: data <= 8'h00;
            16'd8709: data <= 8'hF8;
            16'd8710: data <= 8'h00;
            16'd8711: data <= 8'hF8;
            16'd8712: data <= 8'h00;
            16'd8713: data <= 8'hF8;
            16'd8714: data <= 8'h00;
            16'd8715: data <= 8'hF8;
            16'd8716: data <= 8'h00;
            16'd8717: data <= 8'hF8;
            16'd8718: data <= 8'h00;
            16'd8719: data <= 8'hF8;
            16'd8720: data <= 8'hFF;
            16'd8721: data <= 8'hFF;
            16'd8722: data <= 8'h00;
            16'd8723: data <= 8'hF8;
            16'd8724: data <= 8'h00;
            16'd8725: data <= 8'hF8;
            16'd8726: data <= 8'h00;
            16'd8727: data <= 8'hF8;
            16'd8728: data <= 8'h00;
            16'd8729: data <= 8'hF8;
            16'd8730: data <= 8'h00;
            16'd8731: data <= 8'hF8;
            16'd8732: data <= 8'h00;
            16'd8733: data <= 8'hF8;
            16'd8734: data <= 8'h00;
            16'd8735: data <= 8'hF8;
            16'd8736: data <= 8'h00;
            16'd8737: data <= 8'hF8;
            16'd8738: data <= 8'h00;
            16'd8739: data <= 8'hF8;
            16'd8740: data <= 8'h00;
            16'd8741: data <= 8'hF8;
            16'd8742: data <= 8'h00;
            16'd8743: data <= 8'hF8;
            16'd8744: data <= 8'h00;
            16'd8745: data <= 8'hF8;
            16'd8746: data <= 8'h00;
            16'd8747: data <= 8'hF8;
            16'd8748: data <= 8'h00;
            16'd8749: data <= 8'hF8;
            16'd8750: data <= 8'h00;
            16'd8751: data <= 8'hF8;
            16'd8752: data <= 8'h00;
            16'd8753: data <= 8'hF8;
            16'd8754: data <= 8'h00;
            16'd8755: data <= 8'hF8;
            16'd8756: data <= 8'h00;
            16'd8757: data <= 8'hF8;
            16'd8758: data <= 8'h00;
            16'd8759: data <= 8'hF8;
            16'd8760: data <= 8'hFF;
            16'd8761: data <= 8'hFF;
            16'd8762: data <= 8'h00;
            16'd8763: data <= 8'hF8;
            16'd8764: data <= 8'h00;
            16'd8765: data <= 8'hF8;
            16'd8766: data <= 8'h00;
            16'd8767: data <= 8'hF8;
            16'd8768: data <= 8'h00;
            16'd8769: data <= 8'hF8;
            16'd8770: data <= 8'h00;
            16'd8771: data <= 8'hF8;
            16'd8772: data <= 8'h00;
            16'd8773: data <= 8'hF8;
            16'd8774: data <= 8'h00;
            16'd8775: data <= 8'hF8;
            16'd8776: data <= 8'h00;
            16'd8777: data <= 8'hF8;
            16'd8778: data <= 8'h00;
            16'd8779: data <= 8'hF8;
            16'd8780: data <= 8'h00;
            16'd8781: data <= 8'hF8;
            16'd8782: data <= 8'h00;
            16'd8783: data <= 8'hF8;
            16'd8784: data <= 8'h00;
            16'd8785: data <= 8'hF8;
            16'd8786: data <= 8'h00;
            16'd8787: data <= 8'hF8;
            16'd8788: data <= 8'h00;
            16'd8789: data <= 8'hF8;
            16'd8790: data <= 8'h00;
            16'd8791: data <= 8'hF8;
            16'd8792: data <= 8'h00;
            16'd8793: data <= 8'hF8;
            16'd8794: data <= 8'h00;
            16'd8795: data <= 8'hF8;
            16'd8796: data <= 8'h00;
            16'd8797: data <= 8'hF8;
            16'd8798: data <= 8'h00;
            16'd8799: data <= 8'hF8;
            16'd8800: data <= 8'hFF;
            16'd8801: data <= 8'hFF;
            16'd8802: data <= 8'h00;
            16'd8803: data <= 8'hF8;
            16'd8804: data <= 8'h00;
            16'd8805: data <= 8'hF8;
            16'd8806: data <= 8'h00;
            16'd8807: data <= 8'hF8;
            16'd8808: data <= 8'h00;
            16'd8809: data <= 8'hF8;
            16'd8810: data <= 8'h00;
            16'd8811: data <= 8'hF8;
            16'd8812: data <= 8'h00;
            16'd8813: data <= 8'hF8;
            16'd8814: data <= 8'h00;
            16'd8815: data <= 8'hF8;
            16'd8816: data <= 8'h00;
            16'd8817: data <= 8'hF8;
            16'd8818: data <= 8'h00;
            16'd8819: data <= 8'hF8;
            16'd8820: data <= 8'h00;
            16'd8821: data <= 8'hF8;
            16'd8822: data <= 8'h00;
            16'd8823: data <= 8'hF8;
            16'd8824: data <= 8'h00;
            16'd8825: data <= 8'hF8;
            16'd8826: data <= 8'h00;
            16'd8827: data <= 8'hF8;
            16'd8828: data <= 8'h00;
            16'd8829: data <= 8'hF8;
            16'd8830: data <= 8'h00;
            16'd8831: data <= 8'hF8;
            16'd8832: data <= 8'h00;
            16'd8833: data <= 8'hF8;
            16'd8834: data <= 8'h00;
            16'd8835: data <= 8'hF8;
            16'd8836: data <= 8'h00;
            16'd8837: data <= 8'hF8;
            16'd8838: data <= 8'h00;
            16'd8839: data <= 8'hF8;
            16'd8840: data <= 8'hFF;
            16'd8841: data <= 8'hFF;
            16'd8842: data <= 8'h00;
            16'd8843: data <= 8'hF8;
            16'd8844: data <= 8'h00;
            16'd8845: data <= 8'hF8;
            16'd8846: data <= 8'h00;
            16'd8847: data <= 8'hF8;
            16'd8848: data <= 8'h00;
            16'd8849: data <= 8'hF8;
            16'd8850: data <= 8'h00;
            16'd8851: data <= 8'hF8;
            16'd8852: data <= 8'h00;
            16'd8853: data <= 8'hF8;
            16'd8854: data <= 8'h00;
            16'd8855: data <= 8'hF8;
            16'd8856: data <= 8'h00;
            16'd8857: data <= 8'hF8;
            16'd8858: data <= 8'h00;
            16'd8859: data <= 8'hF8;
            16'd8860: data <= 8'h00;
            16'd8861: data <= 8'hF8;
            16'd8862: data <= 8'h00;
            16'd8863: data <= 8'hF8;
            16'd8864: data <= 8'h00;
            16'd8865: data <= 8'hF8;
            16'd8866: data <= 8'h00;
            16'd8867: data <= 8'hF8;
            16'd8868: data <= 8'h00;
            16'd8869: data <= 8'hF8;
            16'd8870: data <= 8'h00;
            16'd8871: data <= 8'hF8;
            16'd8872: data <= 8'h00;
            16'd8873: data <= 8'hF8;
            16'd8874: data <= 8'h00;
            16'd8875: data <= 8'hF8;
            16'd8876: data <= 8'h00;
            16'd8877: data <= 8'hF8;
            16'd8878: data <= 8'h00;
            16'd8879: data <= 8'hF8;
            16'd8880: data <= 8'hFF;
            16'd8881: data <= 8'hFF;
            16'd8882: data <= 8'h00;
            16'd8883: data <= 8'hF8;
            16'd8884: data <= 8'h00;
            16'd8885: data <= 8'hF8;
            16'd8886: data <= 8'h00;
            16'd8887: data <= 8'hF8;
            16'd8888: data <= 8'h00;
            16'd8889: data <= 8'hF8;
            16'd8890: data <= 8'h00;
            16'd8891: data <= 8'hF8;
            16'd8892: data <= 8'h00;
            16'd8893: data <= 8'hF8;
            16'd8894: data <= 8'h00;
            16'd8895: data <= 8'hF8;
            16'd8896: data <= 8'h00;
            16'd8897: data <= 8'hF8;
            16'd8898: data <= 8'h00;
            16'd8899: data <= 8'hF8;
            16'd8900: data <= 8'h00;
            16'd8901: data <= 8'hF8;
            16'd8902: data <= 8'h00;
            16'd8903: data <= 8'hF8;
            16'd8904: data <= 8'h00;
            16'd8905: data <= 8'hF8;
            16'd8906: data <= 8'h00;
            16'd8907: data <= 8'hF8;
            16'd8908: data <= 8'h00;
            16'd8909: data <= 8'hF8;
            16'd8910: data <= 8'h00;
            16'd8911: data <= 8'hF8;
            16'd8912: data <= 8'h00;
            16'd8913: data <= 8'hF8;
            16'd8914: data <= 8'h00;
            16'd8915: data <= 8'hF8;
            16'd8916: data <= 8'h00;
            16'd8917: data <= 8'hF8;
            16'd8918: data <= 8'h00;
            16'd8919: data <= 8'hF8;
            16'd8920: data <= 8'hFF;
            16'd8921: data <= 8'hFF;
            16'd8922: data <= 8'h00;
            16'd8923: data <= 8'hF8;
            16'd8924: data <= 8'h00;
            16'd8925: data <= 8'hF8;
            16'd8926: data <= 8'h00;
            16'd8927: data <= 8'hF8;
            16'd8928: data <= 8'h00;
            16'd8929: data <= 8'hF8;
            16'd8930: data <= 8'h00;
            16'd8931: data <= 8'hF8;
            16'd8932: data <= 8'h00;
            16'd8933: data <= 8'hF8;
            16'd8934: data <= 8'h00;
            16'd8935: data <= 8'hF8;
            16'd8936: data <= 8'h00;
            16'd8937: data <= 8'hF8;
            16'd8938: data <= 8'h00;
            16'd8939: data <= 8'hF8;
            16'd8940: data <= 8'h00;
            16'd8941: data <= 8'hF8;
            16'd8942: data <= 8'h00;
            16'd8943: data <= 8'hF8;
            16'd8944: data <= 8'h00;
            16'd8945: data <= 8'hF8;
            16'd8946: data <= 8'h00;
            16'd8947: data <= 8'hF8;
            16'd8948: data <= 8'h00;
            16'd8949: data <= 8'hF8;
            16'd8950: data <= 8'h00;
            16'd8951: data <= 8'hF8;
            16'd8952: data <= 8'h00;
            16'd8953: data <= 8'hF8;
            16'd8954: data <= 8'h00;
            16'd8955: data <= 8'hF8;
            16'd8956: data <= 8'h00;
            16'd8957: data <= 8'hF8;
            16'd8958: data <= 8'h00;
            16'd8959: data <= 8'hF8;
            16'd8960: data <= 8'hFF;
            16'd8961: data <= 8'hFF;
            16'd8962: data <= 8'h00;
            16'd8963: data <= 8'hF8;
            16'd8964: data <= 8'h00;
            16'd8965: data <= 8'hF8;
            16'd8966: data <= 8'h00;
            16'd8967: data <= 8'hF8;
            16'd8968: data <= 8'h00;
            16'd8969: data <= 8'hF8;
            16'd8970: data <= 8'h00;
            16'd8971: data <= 8'hF8;
            16'd8972: data <= 8'h00;
            16'd8973: data <= 8'hF8;
            16'd8974: data <= 8'h00;
            16'd8975: data <= 8'hF8;
            16'd8976: data <= 8'h00;
            16'd8977: data <= 8'hF8;
            16'd8978: data <= 8'h00;
            16'd8979: data <= 8'hF8;
            16'd8980: data <= 8'h00;
            16'd8981: data <= 8'hF8;
            16'd8982: data <= 8'h00;
            16'd8983: data <= 8'hF8;
            16'd8984: data <= 8'h00;
            16'd8985: data <= 8'hF8;
            16'd8986: data <= 8'h00;
            16'd8987: data <= 8'hF8;
            16'd8988: data <= 8'h00;
            16'd8989: data <= 8'hF8;
            16'd8990: data <= 8'h00;
            16'd8991: data <= 8'hF8;
            16'd8992: data <= 8'h00;
            16'd8993: data <= 8'hF8;
            16'd8994: data <= 8'h00;
            16'd8995: data <= 8'hF8;
            16'd8996: data <= 8'h00;
            16'd8997: data <= 8'hF8;
            16'd8998: data <= 8'h00;
            16'd8999: data <= 8'hF8;
            16'd9000: data <= 8'hFF;
            16'd9001: data <= 8'hFF;
            16'd9002: data <= 8'h00;
            16'd9003: data <= 8'hF8;
            16'd9004: data <= 8'h00;
            16'd9005: data <= 8'hF8;
            16'd9006: data <= 8'h00;
            16'd9007: data <= 8'hF8;
            16'd9008: data <= 8'h00;
            16'd9009: data <= 8'hF8;
            16'd9010: data <= 8'h00;
            16'd9011: data <= 8'hF8;
            16'd9012: data <= 8'h00;
            16'd9013: data <= 8'hF8;
            16'd9014: data <= 8'h00;
            16'd9015: data <= 8'hF8;
            16'd9016: data <= 8'h00;
            16'd9017: data <= 8'hF8;
            16'd9018: data <= 8'h00;
            16'd9019: data <= 8'hF8;
            16'd9020: data <= 8'h00;
            16'd9021: data <= 8'hF8;
            16'd9022: data <= 8'h00;
            16'd9023: data <= 8'hF8;
            16'd9024: data <= 8'h00;
            16'd9025: data <= 8'hF8;
            16'd9026: data <= 8'h00;
            16'd9027: data <= 8'hF8;
            16'd9028: data <= 8'h00;
            16'd9029: data <= 8'hF8;
            16'd9030: data <= 8'h00;
            16'd9031: data <= 8'hF8;
            16'd9032: data <= 8'h00;
            16'd9033: data <= 8'hF8;
            16'd9034: data <= 8'h00;
            16'd9035: data <= 8'hF8;
            16'd9036: data <= 8'h00;
            16'd9037: data <= 8'hF8;
            16'd9038: data <= 8'h00;
            16'd9039: data <= 8'hF8;
            16'd9040: data <= 8'hFF;
            16'd9041: data <= 8'hFF;
            16'd9042: data <= 8'h00;
            16'd9043: data <= 8'hF8;
            16'd9044: data <= 8'h00;
            16'd9045: data <= 8'hF8;
            16'd9046: data <= 8'h00;
            16'd9047: data <= 8'hF8;
            16'd9048: data <= 8'h00;
            16'd9049: data <= 8'hF8;
            16'd9050: data <= 8'h00;
            16'd9051: data <= 8'hF8;
            16'd9052: data <= 8'h00;
            16'd9053: data <= 8'hF8;
            16'd9054: data <= 8'h00;
            16'd9055: data <= 8'hF8;
            16'd9056: data <= 8'h00;
            16'd9057: data <= 8'hF8;
            16'd9058: data <= 8'h00;
            16'd9059: data <= 8'hF8;
            16'd9060: data <= 8'h00;
            16'd9061: data <= 8'hF8;
            16'd9062: data <= 8'h00;
            16'd9063: data <= 8'hF8;
            16'd9064: data <= 8'h00;
            16'd9065: data <= 8'hF8;
            16'd9066: data <= 8'h00;
            16'd9067: data <= 8'hF8;
            16'd9068: data <= 8'h00;
            16'd9069: data <= 8'hF8;
            16'd9070: data <= 8'h00;
            16'd9071: data <= 8'hF8;
            16'd9072: data <= 8'h00;
            16'd9073: data <= 8'hF8;
            16'd9074: data <= 8'h00;
            16'd9075: data <= 8'hF8;
            16'd9076: data <= 8'h00;
            16'd9077: data <= 8'hF8;
            16'd9078: data <= 8'h00;
            16'd9079: data <= 8'hF8;
            16'd9080: data <= 8'hFF;
            16'd9081: data <= 8'hFF;
            16'd9082: data <= 8'h00;
            16'd9083: data <= 8'hF8;
            16'd9084: data <= 8'h00;
            16'd9085: data <= 8'hF8;
            16'd9086: data <= 8'h00;
            16'd9087: data <= 8'hF8;
            16'd9088: data <= 8'h00;
            16'd9089: data <= 8'hF8;
            16'd9090: data <= 8'h00;
            16'd9091: data <= 8'hF8;
            16'd9092: data <= 8'h00;
            16'd9093: data <= 8'hF8;
            16'd9094: data <= 8'h00;
            16'd9095: data <= 8'hF8;
            16'd9096: data <= 8'h00;
            16'd9097: data <= 8'hF8;
            16'd9098: data <= 8'h00;
            16'd9099: data <= 8'hF8;
            16'd9100: data <= 8'h00;
            16'd9101: data <= 8'hF8;
            16'd9102: data <= 8'h00;
            16'd9103: data <= 8'hF8;
            16'd9104: data <= 8'h00;
            16'd9105: data <= 8'hF8;
            16'd9106: data <= 8'h00;
            16'd9107: data <= 8'hF8;
            16'd9108: data <= 8'h00;
            16'd9109: data <= 8'hF8;
            16'd9110: data <= 8'h00;
            16'd9111: data <= 8'hF8;
            16'd9112: data <= 8'h00;
            16'd9113: data <= 8'hF8;
            16'd9114: data <= 8'h00;
            16'd9115: data <= 8'hF8;
            16'd9116: data <= 8'h00;
            16'd9117: data <= 8'hF8;
            16'd9118: data <= 8'h00;
            16'd9119: data <= 8'hF8;
            16'd9120: data <= 8'hFF;
            16'd9121: data <= 8'hFF;
            16'd9122: data <= 8'h00;
            16'd9123: data <= 8'hF8;
            16'd9124: data <= 8'h00;
            16'd9125: data <= 8'hF8;
            16'd9126: data <= 8'h00;
            16'd9127: data <= 8'hF8;
            16'd9128: data <= 8'h00;
            16'd9129: data <= 8'hF8;
            16'd9130: data <= 8'h00;
            16'd9131: data <= 8'hF8;
            16'd9132: data <= 8'h00;
            16'd9133: data <= 8'hF8;
            16'd9134: data <= 8'h00;
            16'd9135: data <= 8'hF8;
            16'd9136: data <= 8'h00;
            16'd9137: data <= 8'hF8;
            16'd9138: data <= 8'h00;
            16'd9139: data <= 8'hF8;
            16'd9140: data <= 8'h00;
            16'd9141: data <= 8'hF8;
            16'd9142: data <= 8'h00;
            16'd9143: data <= 8'hF8;
            16'd9144: data <= 8'h00;
            16'd9145: data <= 8'hF8;
            16'd9146: data <= 8'h00;
            16'd9147: data <= 8'hF8;
            16'd9148: data <= 8'h00;
            16'd9149: data <= 8'hF8;
            16'd9150: data <= 8'h00;
            16'd9151: data <= 8'hF8;
            16'd9152: data <= 8'h00;
            16'd9153: data <= 8'hF8;
            16'd9154: data <= 8'h00;
            16'd9155: data <= 8'hF8;
            16'd9156: data <= 8'h00;
            16'd9157: data <= 8'hF8;
            16'd9158: data <= 8'h00;
            16'd9159: data <= 8'hF8;
            16'd9160: data <= 8'hFF;
            16'd9161: data <= 8'hFF;
            16'd9162: data <= 8'h00;
            16'd9163: data <= 8'hF8;
            16'd9164: data <= 8'h00;
            16'd9165: data <= 8'hF8;
            16'd9166: data <= 8'h00;
            16'd9167: data <= 8'hF8;
            16'd9168: data <= 8'h00;
            16'd9169: data <= 8'hF8;
            16'd9170: data <= 8'h00;
            16'd9171: data <= 8'hF8;
            16'd9172: data <= 8'h00;
            16'd9173: data <= 8'hF8;
            16'd9174: data <= 8'h00;
            16'd9175: data <= 8'hF8;
            16'd9176: data <= 8'h00;
            16'd9177: data <= 8'hF8;
            16'd9178: data <= 8'h00;
            16'd9179: data <= 8'hF8;
            16'd9180: data <= 8'h00;
            16'd9181: data <= 8'hF8;
            16'd9182: data <= 8'h00;
            16'd9183: data <= 8'hF8;
            16'd9184: data <= 8'h00;
            16'd9185: data <= 8'hF8;
            16'd9186: data <= 8'h00;
            16'd9187: data <= 8'hF8;
            16'd9188: data <= 8'h00;
            16'd9189: data <= 8'hF8;
            16'd9190: data <= 8'h00;
            16'd9191: data <= 8'hF8;
            16'd9192: data <= 8'h00;
            16'd9193: data <= 8'hF8;
            16'd9194: data <= 8'h00;
            16'd9195: data <= 8'hF8;
            16'd9196: data <= 8'h00;
            16'd9197: data <= 8'hF8;
            16'd9198: data <= 8'h00;
            16'd9199: data <= 8'hF8;
            16'd9200: data <= 8'hFF;
            16'd9201: data <= 8'hFF;
            16'd9202: data <= 8'h00;
            16'd9203: data <= 8'hF8;
            16'd9204: data <= 8'h00;
            16'd9205: data <= 8'hF8;
            16'd9206: data <= 8'h00;
            16'd9207: data <= 8'hF8;
            16'd9208: data <= 8'h00;
            16'd9209: data <= 8'hF8;
            16'd9210: data <= 8'h00;
            16'd9211: data <= 8'hF8;
            16'd9212: data <= 8'h00;
            16'd9213: data <= 8'hF8;
            16'd9214: data <= 8'h00;
            16'd9215: data <= 8'hF8;
            16'd9216: data <= 8'h00;
            16'd9217: data <= 8'hF8;
            16'd9218: data <= 8'h00;
            16'd9219: data <= 8'hF8;
            16'd9220: data <= 8'h00;
            16'd9221: data <= 8'hF8;
            16'd9222: data <= 8'h00;
            16'd9223: data <= 8'hF8;
            16'd9224: data <= 8'h00;
            16'd9225: data <= 8'hF8;
            16'd9226: data <= 8'h00;
            16'd9227: data <= 8'hF8;
            16'd9228: data <= 8'h00;
            16'd9229: data <= 8'hF8;
            16'd9230: data <= 8'h00;
            16'd9231: data <= 8'hF8;
            16'd9232: data <= 8'h00;
            16'd9233: data <= 8'hF8;
            16'd9234: data <= 8'h00;
            16'd9235: data <= 8'hF8;
            16'd9236: data <= 8'h00;
            16'd9237: data <= 8'hF8;
            16'd9238: data <= 8'h00;
            16'd9239: data <= 8'hF8;
            16'd9240: data <= 8'hFF;
            16'd9241: data <= 8'hFF;
            16'd9242: data <= 8'h00;
            16'd9243: data <= 8'hF8;
            16'd9244: data <= 8'h00;
            16'd9245: data <= 8'hF8;
            16'd9246: data <= 8'h00;
            16'd9247: data <= 8'hF8;
            16'd9248: data <= 8'h00;
            16'd9249: data <= 8'hF8;
            16'd9250: data <= 8'h00;
            16'd9251: data <= 8'hF8;
            16'd9252: data <= 8'h00;
            16'd9253: data <= 8'hF8;
            16'd9254: data <= 8'h00;
            16'd9255: data <= 8'hF8;
            16'd9256: data <= 8'h00;
            16'd9257: data <= 8'hF8;
            16'd9258: data <= 8'h00;
            16'd9259: data <= 8'hF8;
            16'd9260: data <= 8'h00;
            16'd9261: data <= 8'hF8;
            16'd9262: data <= 8'h00;
            16'd9263: data <= 8'hF8;
            16'd9264: data <= 8'h00;
            16'd9265: data <= 8'hF8;
            16'd9266: data <= 8'h00;
            16'd9267: data <= 8'hF8;
            16'd9268: data <= 8'h00;
            16'd9269: data <= 8'hF8;
            16'd9270: data <= 8'h00;
            16'd9271: data <= 8'hF8;
            16'd9272: data <= 8'h00;
            16'd9273: data <= 8'hF8;
            16'd9274: data <= 8'h00;
            16'd9275: data <= 8'hF8;
            16'd9276: data <= 8'h00;
            16'd9277: data <= 8'hF8;
            16'd9278: data <= 8'h00;
            16'd9279: data <= 8'hF8;
            16'd9280: data <= 8'hFF;
            16'd9281: data <= 8'hFF;
            16'd9282: data <= 8'h00;
            16'd9283: data <= 8'hF8;
            16'd9284: data <= 8'h00;
            16'd9285: data <= 8'hF8;
            16'd9286: data <= 8'h00;
            16'd9287: data <= 8'hF8;
            16'd9288: data <= 8'h00;
            16'd9289: data <= 8'hF8;
            16'd9290: data <= 8'h00;
            16'd9291: data <= 8'hF8;
            16'd9292: data <= 8'h00;
            16'd9293: data <= 8'hF8;
            16'd9294: data <= 8'h00;
            16'd9295: data <= 8'hF8;
            16'd9296: data <= 8'h00;
            16'd9297: data <= 8'hF8;
            16'd9298: data <= 8'h00;
            16'd9299: data <= 8'hF8;
            16'd9300: data <= 8'h00;
            16'd9301: data <= 8'hF8;
            16'd9302: data <= 8'h00;
            16'd9303: data <= 8'hF8;
            16'd9304: data <= 8'h00;
            16'd9305: data <= 8'hF8;
            16'd9306: data <= 8'h00;
            16'd9307: data <= 8'hF8;
            16'd9308: data <= 8'h00;
            16'd9309: data <= 8'hF8;
            16'd9310: data <= 8'h00;
            16'd9311: data <= 8'hF8;
            16'd9312: data <= 8'h00;
            16'd9313: data <= 8'hF8;
            16'd9314: data <= 8'h00;
            16'd9315: data <= 8'hF8;
            16'd9316: data <= 8'h00;
            16'd9317: data <= 8'hF8;
            16'd9318: data <= 8'h00;
            16'd9319: data <= 8'hF8;
            16'd9320: data <= 8'hFF;
            16'd9321: data <= 8'hFF;
            16'd9322: data <= 8'h00;
            16'd9323: data <= 8'hF8;
            16'd9324: data <= 8'h00;
            16'd9325: data <= 8'hF8;
            16'd9326: data <= 8'h00;
            16'd9327: data <= 8'hF8;
            16'd9328: data <= 8'h00;
            16'd9329: data <= 8'hF8;
            16'd9330: data <= 8'h00;
            16'd9331: data <= 8'hF8;
            16'd9332: data <= 8'h00;
            16'd9333: data <= 8'hF8;
            16'd9334: data <= 8'h00;
            16'd9335: data <= 8'hF8;
            16'd9336: data <= 8'h00;
            16'd9337: data <= 8'hF8;
            16'd9338: data <= 8'h00;
            16'd9339: data <= 8'hF8;
            16'd9340: data <= 8'h00;
            16'd9341: data <= 8'hF8;
            16'd9342: data <= 8'h00;
            16'd9343: data <= 8'hF8;
            16'd9344: data <= 8'h00;
            16'd9345: data <= 8'hF8;
            16'd9346: data <= 8'h00;
            16'd9347: data <= 8'hF8;
            16'd9348: data <= 8'h00;
            16'd9349: data <= 8'hF8;
            16'd9350: data <= 8'h00;
            16'd9351: data <= 8'hF8;
            16'd9352: data <= 8'h00;
            16'd9353: data <= 8'hF8;
            16'd9354: data <= 8'h00;
            16'd9355: data <= 8'hF8;
            16'd9356: data <= 8'h00;
            16'd9357: data <= 8'hF8;
            16'd9358: data <= 8'h00;
            16'd9359: data <= 8'hF8;
            16'd9360: data <= 8'hFF;
            16'd9361: data <= 8'hFF;
            16'd9362: data <= 8'h00;
            16'd9363: data <= 8'hF8;
            16'd9364: data <= 8'h00;
            16'd9365: data <= 8'hF8;
            16'd9366: data <= 8'h00;
            16'd9367: data <= 8'hF8;
            16'd9368: data <= 8'h00;
            16'd9369: data <= 8'hF8;
            16'd9370: data <= 8'h00;
            16'd9371: data <= 8'hF8;
            16'd9372: data <= 8'h00;
            16'd9373: data <= 8'hF8;
            16'd9374: data <= 8'h00;
            16'd9375: data <= 8'hF8;
            16'd9376: data <= 8'h00;
            16'd9377: data <= 8'hF8;
            16'd9378: data <= 8'h00;
            16'd9379: data <= 8'hF8;
            16'd9380: data <= 8'h00;
            16'd9381: data <= 8'hF8;
            16'd9382: data <= 8'h00;
            16'd9383: data <= 8'hF8;
            16'd9384: data <= 8'h00;
            16'd9385: data <= 8'hF8;
            16'd9386: data <= 8'h00;
            16'd9387: data <= 8'hF8;
            16'd9388: data <= 8'h00;
            16'd9389: data <= 8'hF8;
            16'd9390: data <= 8'h00;
            16'd9391: data <= 8'hF8;
            16'd9392: data <= 8'h00;
            16'd9393: data <= 8'hF8;
            16'd9394: data <= 8'h00;
            16'd9395: data <= 8'hF8;
            16'd9396: data <= 8'h00;
            16'd9397: data <= 8'hF8;
            16'd9398: data <= 8'h00;
            16'd9399: data <= 8'hF8;
            16'd9400: data <= 8'hFF;
            16'd9401: data <= 8'hFF;
            16'd9402: data <= 8'h00;
            16'd9403: data <= 8'hF8;
            16'd9404: data <= 8'h00;
            16'd9405: data <= 8'hF8;
            16'd9406: data <= 8'h00;
            16'd9407: data <= 8'hF8;
            16'd9408: data <= 8'h00;
            16'd9409: data <= 8'hF8;
            16'd9410: data <= 8'h00;
            16'd9411: data <= 8'hF8;
            16'd9412: data <= 8'h00;
            16'd9413: data <= 8'hF8;
            16'd9414: data <= 8'h00;
            16'd9415: data <= 8'hF8;
            16'd9416: data <= 8'h00;
            16'd9417: data <= 8'hF8;
            16'd9418: data <= 8'h00;
            16'd9419: data <= 8'hF8;
            16'd9420: data <= 8'h00;
            16'd9421: data <= 8'hF8;
            16'd9422: data <= 8'h00;
            16'd9423: data <= 8'hF8;
            16'd9424: data <= 8'h00;
            16'd9425: data <= 8'hF8;
            16'd9426: data <= 8'h00;
            16'd9427: data <= 8'hF8;
            16'd9428: data <= 8'h00;
            16'd9429: data <= 8'hF8;
            16'd9430: data <= 8'h00;
            16'd9431: data <= 8'hF8;
            16'd9432: data <= 8'h00;
            16'd9433: data <= 8'hF8;
            16'd9434: data <= 8'h00;
            16'd9435: data <= 8'hF8;
            16'd9436: data <= 8'h00;
            16'd9437: data <= 8'hF8;
            16'd9438: data <= 8'h00;
            16'd9439: data <= 8'hF8;
            16'd9440: data <= 8'hFF;
            16'd9441: data <= 8'hFF;
            16'd9442: data <= 8'h00;
            16'd9443: data <= 8'hF8;
            16'd9444: data <= 8'h00;
            16'd9445: data <= 8'hF8;
            16'd9446: data <= 8'h00;
            16'd9447: data <= 8'hF8;
            16'd9448: data <= 8'h00;
            16'd9449: data <= 8'hF8;
            16'd9450: data <= 8'h00;
            16'd9451: data <= 8'hF8;
            16'd9452: data <= 8'h00;
            16'd9453: data <= 8'hF8;
            16'd9454: data <= 8'h00;
            16'd9455: data <= 8'hF8;
            16'd9456: data <= 8'h00;
            16'd9457: data <= 8'hF8;
            16'd9458: data <= 8'h00;
            16'd9459: data <= 8'hF8;
            16'd9460: data <= 8'h00;
            16'd9461: data <= 8'hF8;
            16'd9462: data <= 8'h00;
            16'd9463: data <= 8'hF8;
            16'd9464: data <= 8'h00;
            16'd9465: data <= 8'hF8;
            16'd9466: data <= 8'h00;
            16'd9467: data <= 8'hF8;
            16'd9468: data <= 8'h00;
            16'd9469: data <= 8'hF8;
            16'd9470: data <= 8'h00;
            16'd9471: data <= 8'hF8;
            16'd9472: data <= 8'h00;
            16'd9473: data <= 8'hF8;
            16'd9474: data <= 8'h00;
            16'd9475: data <= 8'hF8;
            16'd9476: data <= 8'h00;
            16'd9477: data <= 8'hF8;
            16'd9478: data <= 8'h00;
            16'd9479: data <= 8'hF8;
            16'd9480: data <= 8'hFF;
            16'd9481: data <= 8'hFF;
            16'd9482: data <= 8'h00;
            16'd9483: data <= 8'hF8;
            16'd9484: data <= 8'h00;
            16'd9485: data <= 8'hF8;
            16'd9486: data <= 8'h00;
            16'd9487: data <= 8'hF8;
            16'd9488: data <= 8'h00;
            16'd9489: data <= 8'hF8;
            16'd9490: data <= 8'h00;
            16'd9491: data <= 8'hF8;
            16'd9492: data <= 8'h00;
            16'd9493: data <= 8'hF8;
            16'd9494: data <= 8'h00;
            16'd9495: data <= 8'hF8;
            16'd9496: data <= 8'h00;
            16'd9497: data <= 8'hF8;
            16'd9498: data <= 8'h00;
            16'd9499: data <= 8'hF8;
            16'd9500: data <= 8'h00;
            16'd9501: data <= 8'hF8;
            16'd9502: data <= 8'h00;
            16'd9503: data <= 8'hF8;
            16'd9504: data <= 8'h00;
            16'd9505: data <= 8'hF8;
            16'd9506: data <= 8'h00;
            16'd9507: data <= 8'hF8;
            16'd9508: data <= 8'h00;
            16'd9509: data <= 8'hF8;
            16'd9510: data <= 8'h00;
            16'd9511: data <= 8'hF8;
            16'd9512: data <= 8'h00;
            16'd9513: data <= 8'hF8;
            16'd9514: data <= 8'h00;
            16'd9515: data <= 8'hF8;
            16'd9516: data <= 8'h00;
            16'd9517: data <= 8'hF8;
            16'd9518: data <= 8'h00;
            16'd9519: data <= 8'hF8;
            16'd9520: data <= 8'hFF;
            16'd9521: data <= 8'hFF;
            16'd9522: data <= 8'h00;
            16'd9523: data <= 8'hF8;
            16'd9524: data <= 8'h00;
            16'd9525: data <= 8'hF8;
            16'd9526: data <= 8'h00;
            16'd9527: data <= 8'hF8;
            16'd9528: data <= 8'h00;
            16'd9529: data <= 8'hF8;
            16'd9530: data <= 8'h00;
            16'd9531: data <= 8'hF8;
            16'd9532: data <= 8'h00;
            16'd9533: data <= 8'hF8;
            16'd9534: data <= 8'h00;
            16'd9535: data <= 8'hF8;
            16'd9536: data <= 8'h00;
            16'd9537: data <= 8'hF8;
            16'd9538: data <= 8'h00;
            16'd9539: data <= 8'hF8;
            16'd9540: data <= 8'h00;
            16'd9541: data <= 8'hF8;
            16'd9542: data <= 8'h00;
            16'd9543: data <= 8'hF8;
            16'd9544: data <= 8'h00;
            16'd9545: data <= 8'hF8;
            16'd9546: data <= 8'h00;
            16'd9547: data <= 8'hF8;
            16'd9548: data <= 8'h00;
            16'd9549: data <= 8'hF8;
            16'd9550: data <= 8'h00;
            16'd9551: data <= 8'hF8;
            16'd9552: data <= 8'h00;
            16'd9553: data <= 8'hF8;
            16'd9554: data <= 8'h00;
            16'd9555: data <= 8'hF8;
            16'd9556: data <= 8'h00;
            16'd9557: data <= 8'hF8;
            16'd9558: data <= 8'h00;
            16'd9559: data <= 8'hF8;
            16'd9560: data <= 8'hFF;
            16'd9561: data <= 8'hFF;
            16'd9562: data <= 8'h00;
            16'd9563: data <= 8'hF8;
            16'd9564: data <= 8'h00;
            16'd9565: data <= 8'hF8;
            16'd9566: data <= 8'h00;
            16'd9567: data <= 8'hF8;
            16'd9568: data <= 8'h00;
            16'd9569: data <= 8'hF8;
            16'd9570: data <= 8'h00;
            16'd9571: data <= 8'hF8;
            16'd9572: data <= 8'h00;
            16'd9573: data <= 8'hF8;
            16'd9574: data <= 8'h00;
            16'd9575: data <= 8'hF8;
            16'd9576: data <= 8'h00;
            16'd9577: data <= 8'hF8;
            16'd9578: data <= 8'h00;
            16'd9579: data <= 8'hF8;
            16'd9580: data <= 8'h00;
            16'd9581: data <= 8'hF8;
            16'd9582: data <= 8'h00;
            16'd9583: data <= 8'hF8;
            16'd9584: data <= 8'h00;
            16'd9585: data <= 8'hF8;
            16'd9586: data <= 8'h00;
            16'd9587: data <= 8'hF8;
            16'd9588: data <= 8'h00;
            16'd9589: data <= 8'hF8;
            16'd9590: data <= 8'h00;
            16'd9591: data <= 8'hF8;
            16'd9592: data <= 8'h00;
            16'd9593: data <= 8'hF8;
            16'd9594: data <= 8'h00;
            16'd9595: data <= 8'hF8;
            16'd9596: data <= 8'h00;
            16'd9597: data <= 8'hF8;
            16'd9598: data <= 8'h00;
            16'd9599: data <= 8'hF8;
            16'd9600: data <= 8'hFF;
            16'd9601: data <= 8'hFF;
            16'd9602: data <= 8'hFF;
            16'd9603: data <= 8'hFF;
            16'd9604: data <= 8'hFF;
            16'd9605: data <= 8'hFF;
            16'd9606: data <= 8'hFF;
            16'd9607: data <= 8'hFF;
            16'd9608: data <= 8'hFF;
            16'd9609: data <= 8'hFF;
            16'd9610: data <= 8'hFF;
            16'd9611: data <= 8'hFF;
            16'd9612: data <= 8'hFF;
            16'd9613: data <= 8'hFF;
            16'd9614: data <= 8'hFF;
            16'd9615: data <= 8'hFF;
            16'd9616: data <= 8'hFF;
            16'd9617: data <= 8'hFF;
            16'd9618: data <= 8'hFF;
            16'd9619: data <= 8'hFF;
            16'd9620: data <= 8'hFF;
            16'd9621: data <= 8'hFF;
            16'd9622: data <= 8'hFF;
            16'd9623: data <= 8'hFF;
            16'd9624: data <= 8'hFF;
            16'd9625: data <= 8'hFF;
            16'd9626: data <= 8'hFF;
            16'd9627: data <= 8'hFF;
            16'd9628: data <= 8'hFF;
            16'd9629: data <= 8'hFF;
            16'd9630: data <= 8'hFF;
            16'd9631: data <= 8'hFF;
            16'd9632: data <= 8'hFF;
            16'd9633: data <= 8'hFF;
            16'd9634: data <= 8'hFF;
            16'd9635: data <= 8'hFF;
            16'd9636: data <= 8'hFF;
            16'd9637: data <= 8'hFF;
            16'd9638: data <= 8'hFF;
            16'd9639: data <= 8'hFF;
            16'd9640: data <= 8'hFF;
            16'd9641: data <= 8'hFF;
            16'd9642: data <= 8'hFF;
            16'd9643: data <= 8'hFF;
            16'd9644: data <= 8'hFF;
            16'd9645: data <= 8'hFF;
            16'd9646: data <= 8'hFF;
            16'd9647: data <= 8'hFF;
            16'd9648: data <= 8'hFF;
            16'd9649: data <= 8'hFF;
            16'd9650: data <= 8'hFF;
            16'd9651: data <= 8'hFF;
            16'd9652: data <= 8'hFF;
            16'd9653: data <= 8'hFF;
            16'd9654: data <= 8'hFF;
            16'd9655: data <= 8'hFF;
            16'd9656: data <= 8'hFF;
            16'd9657: data <= 8'hFF;
            16'd9658: data <= 8'hFF;
            16'd9659: data <= 8'hFF;
            16'd9660: data <= 8'hFF;
            16'd9661: data <= 8'hFF;
            16'd9662: data <= 8'hFF;
            16'd9663: data <= 8'hFF;
            16'd9664: data <= 8'hFF;
            16'd9665: data <= 8'hFF;
            16'd9666: data <= 8'hFF;
            16'd9667: data <= 8'hFF;
            16'd9668: data <= 8'hFF;
            16'd9669: data <= 8'hFF;
            16'd9670: data <= 8'hFF;
            16'd9671: data <= 8'hFF;
            16'd9672: data <= 8'hFF;
            16'd9673: data <= 8'hFF;
            16'd9674: data <= 8'hFF;
            16'd9675: data <= 8'hFF;
            16'd9676: data <= 8'hFF;
            16'd9677: data <= 8'hFF;
            16'd9678: data <= 8'hFF;
            16'd9679: data <= 8'hFF;
            16'd9680: data <= 8'hFF;
            16'd9681: data <= 8'hFF;
            16'd9682: data <= 8'hFF;
            16'd9683: data <= 8'hFF;
            16'd9684: data <= 8'hFF;
            16'd9685: data <= 8'hFF;
            16'd9686: data <= 8'hFF;
            16'd9687: data <= 8'hFF;
            16'd9688: data <= 8'hFF;
            16'd9689: data <= 8'hFF;
            16'd9690: data <= 8'hFF;
            16'd9691: data <= 8'hFF;
            16'd9692: data <= 8'hFF;
            16'd9693: data <= 8'hFF;
            16'd9694: data <= 8'hFF;
            16'd9695: data <= 8'hFF;
            16'd9696: data <= 8'hFF;
            16'd9697: data <= 8'hFF;
            16'd9698: data <= 8'hFF;
            16'd9699: data <= 8'hFF;
            16'd9700: data <= 8'hFF;
            16'd9701: data <= 8'hFF;
            16'd9702: data <= 8'hFF;
            16'd9703: data <= 8'hFF;
            16'd9704: data <= 8'hFF;
            16'd9705: data <= 8'hFF;
            16'd9706: data <= 8'hFF;
            16'd9707: data <= 8'hFF;
            16'd9708: data <= 8'hFF;
            16'd9709: data <= 8'hFF;
            16'd9710: data <= 8'hFF;
            16'd9711: data <= 8'hFF;
            16'd9712: data <= 8'hFF;
            16'd9713: data <= 8'hFF;
            16'd9714: data <= 8'hFF;
            16'd9715: data <= 8'hFF;
            16'd9716: data <= 8'hFF;
            16'd9717: data <= 8'hFF;
            16'd9718: data <= 8'hFF;
            16'd9719: data <= 8'hFF;
            16'd9720: data <= 8'hFF;
            16'd9721: data <= 8'hFF;
            16'd9722: data <= 8'hFF;
            16'd9723: data <= 8'hFF;
            16'd9724: data <= 8'hFF;
            16'd9725: data <= 8'hFF;
            16'd9726: data <= 8'hFF;
            16'd9727: data <= 8'hFF;
            16'd9728: data <= 8'hFF;
            16'd9729: data <= 8'hFF;
            16'd9730: data <= 8'hFF;
            16'd9731: data <= 8'hFF;
            16'd9732: data <= 8'hFF;
            16'd9733: data <= 8'hFF;
            16'd9734: data <= 8'hFF;
            16'd9735: data <= 8'hFF;
            16'd9736: data <= 8'hFF;
            16'd9737: data <= 8'hFF;
            16'd9738: data <= 8'hFF;
            16'd9739: data <= 8'hFF;
            16'd9740: data <= 8'hFF;
            16'd9741: data <= 8'hFF;
            16'd9742: data <= 8'hFF;
            16'd9743: data <= 8'hFF;
            16'd9744: data <= 8'hFF;
            16'd9745: data <= 8'hFF;
            16'd9746: data <= 8'hFF;
            16'd9747: data <= 8'hFF;
            16'd9748: data <= 8'hFF;
            16'd9749: data <= 8'hFF;
            16'd9750: data <= 8'hFF;
            16'd9751: data <= 8'hFF;
            16'd9752: data <= 8'hFF;
            16'd9753: data <= 8'hFF;
            16'd9754: data <= 8'hFF;
            16'd9755: data <= 8'hFF;
            16'd9756: data <= 8'hFF;
            16'd9757: data <= 8'hFF;
            16'd9758: data <= 8'hFF;
            16'd9759: data <= 8'hFF;
            16'd9760: data <= 8'hFF;
            16'd9761: data <= 8'hFF;
            16'd9762: data <= 8'hFF;
            16'd9763: data <= 8'hFF;
            16'd9764: data <= 8'hFF;
            16'd9765: data <= 8'hFF;
            16'd9766: data <= 8'hFF;
            16'd9767: data <= 8'hFF;
            16'd9768: data <= 8'hFF;
            16'd9769: data <= 8'hFF;
            16'd9770: data <= 8'hFF;
            16'd9771: data <= 8'hFF;
            16'd9772: data <= 8'hFF;
            16'd9773: data <= 8'hFF;
            16'd9774: data <= 8'hFF;
            16'd9775: data <= 8'hFF;
            16'd9776: data <= 8'hFF;
            16'd9777: data <= 8'hFF;
            16'd9778: data <= 8'hFF;
            16'd9779: data <= 8'hFF;
            16'd9780: data <= 8'hFF;
            16'd9781: data <= 8'hFF;
            16'd9782: data <= 8'hFF;
            16'd9783: data <= 8'hFF;
            16'd9784: data <= 8'hFF;
            16'd9785: data <= 8'hFF;
            16'd9786: data <= 8'hFF;
            16'd9787: data <= 8'hFF;
            16'd9788: data <= 8'hFF;
            16'd9789: data <= 8'hFF;
            16'd9790: data <= 8'hFF;
            16'd9791: data <= 8'hFF;
            16'd9792: data <= 8'hFF;
            16'd9793: data <= 8'hFF;
            16'd9794: data <= 8'hFF;
            16'd9795: data <= 8'hFF;
            16'd9796: data <= 8'hFF;
            16'd9797: data <= 8'hFF;
            16'd9798: data <= 8'hFF;
            16'd9799: data <= 8'hFF;
            16'd9800: data <= 8'hFF;
            16'd9801: data <= 8'hFF;
            16'd9802: data <= 8'hFF;
            16'd9803: data <= 8'hFF;
            16'd9804: data <= 8'hFF;
            16'd9805: data <= 8'hFF;
            16'd9806: data <= 8'hFF;
            16'd9807: data <= 8'hFF;
            16'd9808: data <= 8'hFF;
            16'd9809: data <= 8'hFF;
            16'd9810: data <= 8'hFF;
            16'd9811: data <= 8'hFF;
            16'd9812: data <= 8'hFF;
            16'd9813: data <= 8'hFF;
            16'd9814: data <= 8'hFF;
            16'd9815: data <= 8'hFF;
            16'd9816: data <= 8'hFF;
            16'd9817: data <= 8'hFF;
            16'd9818: data <= 8'hFF;
            16'd9819: data <= 8'hFF;
            16'd9820: data <= 8'hFF;
            16'd9821: data <= 8'hFF;
            16'd9822: data <= 8'hFF;
            16'd9823: data <= 8'hFF;
            16'd9824: data <= 8'hFF;
            16'd9825: data <= 8'hFF;
            16'd9826: data <= 8'hFF;
            16'd9827: data <= 8'hFF;
            16'd9828: data <= 8'hFF;
            16'd9829: data <= 8'hFF;
            16'd9830: data <= 8'hFF;
            16'd9831: data <= 8'hFF;
            16'd9832: data <= 8'hFF;
            16'd9833: data <= 8'hFF;
            16'd9834: data <= 8'hFF;
            16'd9835: data <= 8'hFF;
            16'd9836: data <= 8'hFF;
            16'd9837: data <= 8'hFF;
            16'd9838: data <= 8'hFF;
            16'd9839: data <= 8'hFF;
            16'd9840: data <= 8'hFF;
            16'd9841: data <= 8'hFF;
            16'd9842: data <= 8'h00;
            16'd9843: data <= 8'hF8;
            16'd9844: data <= 8'h00;
            16'd9845: data <= 8'hF8;
            16'd9846: data <= 8'h00;
            16'd9847: data <= 8'hF8;
            16'd9848: data <= 8'h00;
            16'd9849: data <= 8'hF8;
            16'd9850: data <= 8'h00;
            16'd9851: data <= 8'hF8;
            16'd9852: data <= 8'h00;
            16'd9853: data <= 8'hF8;
            16'd9854: data <= 8'h00;
            16'd9855: data <= 8'hF8;
            16'd9856: data <= 8'h00;
            16'd9857: data <= 8'hF8;
            16'd9858: data <= 8'h00;
            16'd9859: data <= 8'hF8;
            16'd9860: data <= 8'h00;
            16'd9861: data <= 8'hF8;
            16'd9862: data <= 8'h00;
            16'd9863: data <= 8'hF8;
            16'd9864: data <= 8'h00;
            16'd9865: data <= 8'hF8;
            16'd9866: data <= 8'h00;
            16'd9867: data <= 8'hF8;
            16'd9868: data <= 8'h00;
            16'd9869: data <= 8'hF8;
            16'd9870: data <= 8'h00;
            16'd9871: data <= 8'hF8;
            16'd9872: data <= 8'h00;
            16'd9873: data <= 8'hF8;
            16'd9874: data <= 8'h00;
            16'd9875: data <= 8'hF8;
            16'd9876: data <= 8'h00;
            16'd9877: data <= 8'hF8;
            16'd9878: data <= 8'h00;
            16'd9879: data <= 8'hF8;
            16'd9880: data <= 8'hFF;
            16'd9881: data <= 8'hFF;
            16'd9882: data <= 8'h00;
            16'd9883: data <= 8'hF8;
            16'd9884: data <= 8'h00;
            16'd9885: data <= 8'hF8;
            16'd9886: data <= 8'h00;
            16'd9887: data <= 8'hF8;
            16'd9888: data <= 8'h00;
            16'd9889: data <= 8'hF8;
            16'd9890: data <= 8'h00;
            16'd9891: data <= 8'hF8;
            16'd9892: data <= 8'h00;
            16'd9893: data <= 8'hF8;
            16'd9894: data <= 8'h00;
            16'd9895: data <= 8'hF8;
            16'd9896: data <= 8'h00;
            16'd9897: data <= 8'hF8;
            16'd9898: data <= 8'h00;
            16'd9899: data <= 8'hF8;
            16'd9900: data <= 8'h00;
            16'd9901: data <= 8'hF8;
            16'd9902: data <= 8'h00;
            16'd9903: data <= 8'hF8;
            16'd9904: data <= 8'h00;
            16'd9905: data <= 8'hF8;
            16'd9906: data <= 8'h00;
            16'd9907: data <= 8'hF8;
            16'd9908: data <= 8'h00;
            16'd9909: data <= 8'hF8;
            16'd9910: data <= 8'h00;
            16'd9911: data <= 8'hF8;
            16'd9912: data <= 8'h00;
            16'd9913: data <= 8'hF8;
            16'd9914: data <= 8'h00;
            16'd9915: data <= 8'hF8;
            16'd9916: data <= 8'h00;
            16'd9917: data <= 8'hF8;
            16'd9918: data <= 8'h00;
            16'd9919: data <= 8'hF8;
            16'd9920: data <= 8'hFF;
            16'd9921: data <= 8'hFF;
            16'd9922: data <= 8'h00;
            16'd9923: data <= 8'hF8;
            16'd9924: data <= 8'h00;
            16'd9925: data <= 8'hF8;
            16'd9926: data <= 8'h00;
            16'd9927: data <= 8'hF8;
            16'd9928: data <= 8'h00;
            16'd9929: data <= 8'hF8;
            16'd9930: data <= 8'h00;
            16'd9931: data <= 8'hF8;
            16'd9932: data <= 8'h00;
            16'd9933: data <= 8'hF8;
            16'd9934: data <= 8'h00;
            16'd9935: data <= 8'hF8;
            16'd9936: data <= 8'h00;
            16'd9937: data <= 8'hF8;
            16'd9938: data <= 8'h00;
            16'd9939: data <= 8'hF8;
            16'd9940: data <= 8'h00;
            16'd9941: data <= 8'hF8;
            16'd9942: data <= 8'h00;
            16'd9943: data <= 8'hF8;
            16'd9944: data <= 8'h00;
            16'd9945: data <= 8'hF8;
            16'd9946: data <= 8'h00;
            16'd9947: data <= 8'hF8;
            16'd9948: data <= 8'h00;
            16'd9949: data <= 8'hF8;
            16'd9950: data <= 8'h00;
            16'd9951: data <= 8'hF8;
            16'd9952: data <= 8'h00;
            16'd9953: data <= 8'hF8;
            16'd9954: data <= 8'h00;
            16'd9955: data <= 8'hF8;
            16'd9956: data <= 8'h00;
            16'd9957: data <= 8'hF8;
            16'd9958: data <= 8'h00;
            16'd9959: data <= 8'hF8;
            16'd9960: data <= 8'hFF;
            16'd9961: data <= 8'hFF;
            16'd9962: data <= 8'h00;
            16'd9963: data <= 8'hF8;
            16'd9964: data <= 8'h00;
            16'd9965: data <= 8'hF8;
            16'd9966: data <= 8'h00;
            16'd9967: data <= 8'hF8;
            16'd9968: data <= 8'h00;
            16'd9969: data <= 8'hF8;
            16'd9970: data <= 8'h00;
            16'd9971: data <= 8'hF8;
            16'd9972: data <= 8'h00;
            16'd9973: data <= 8'hF8;
            16'd9974: data <= 8'h00;
            16'd9975: data <= 8'hF8;
            16'd9976: data <= 8'h00;
            16'd9977: data <= 8'hF8;
            16'd9978: data <= 8'h00;
            16'd9979: data <= 8'hF8;
            16'd9980: data <= 8'h00;
            16'd9981: data <= 8'hF8;
            16'd9982: data <= 8'h00;
            16'd9983: data <= 8'hF8;
            16'd9984: data <= 8'h00;
            16'd9985: data <= 8'hF8;
            16'd9986: data <= 8'h00;
            16'd9987: data <= 8'hF8;
            16'd9988: data <= 8'h00;
            16'd9989: data <= 8'hF8;
            16'd9990: data <= 8'h00;
            16'd9991: data <= 8'hF8;
            16'd9992: data <= 8'h00;
            16'd9993: data <= 8'hF8;
            16'd9994: data <= 8'h00;
            16'd9995: data <= 8'hF8;
            16'd9996: data <= 8'h00;
            16'd9997: data <= 8'hF8;
            16'd9998: data <= 8'h00;
            16'd9999: data <= 8'hF8;
            16'd10000: data <= 8'hFF;
            16'd10001: data <= 8'hFF;
            16'd10002: data <= 8'h00;
            16'd10003: data <= 8'hF8;
            16'd10004: data <= 8'h00;
            16'd10005: data <= 8'hF8;
            16'd10006: data <= 8'h00;
            16'd10007: data <= 8'hF8;
            16'd10008: data <= 8'h00;
            16'd10009: data <= 8'hF8;
            16'd10010: data <= 8'h00;
            16'd10011: data <= 8'hF8;
            16'd10012: data <= 8'h00;
            16'd10013: data <= 8'hF8;
            16'd10014: data <= 8'h00;
            16'd10015: data <= 8'hF8;
            16'd10016: data <= 8'h00;
            16'd10017: data <= 8'hF8;
            16'd10018: data <= 8'h00;
            16'd10019: data <= 8'hF8;
            16'd10020: data <= 8'h00;
            16'd10021: data <= 8'hF8;
            16'd10022: data <= 8'h00;
            16'd10023: data <= 8'hF8;
            16'd10024: data <= 8'h00;
            16'd10025: data <= 8'hF8;
            16'd10026: data <= 8'h00;
            16'd10027: data <= 8'hF8;
            16'd10028: data <= 8'h00;
            16'd10029: data <= 8'hF8;
            16'd10030: data <= 8'h00;
            16'd10031: data <= 8'hF8;
            16'd10032: data <= 8'h00;
            16'd10033: data <= 8'hF8;
            16'd10034: data <= 8'h00;
            16'd10035: data <= 8'hF8;
            16'd10036: data <= 8'h00;
            16'd10037: data <= 8'hF8;
            16'd10038: data <= 8'h00;
            16'd10039: data <= 8'hF8;
            16'd10040: data <= 8'hFF;
            16'd10041: data <= 8'hFF;
            16'd10042: data <= 8'h00;
            16'd10043: data <= 8'hF8;
            16'd10044: data <= 8'h00;
            16'd10045: data <= 8'hF8;
            16'd10046: data <= 8'h00;
            16'd10047: data <= 8'hF8;
            16'd10048: data <= 8'h00;
            16'd10049: data <= 8'hF8;
            16'd10050: data <= 8'h00;
            16'd10051: data <= 8'hF8;
            16'd10052: data <= 8'h00;
            16'd10053: data <= 8'hF8;
            16'd10054: data <= 8'h00;
            16'd10055: data <= 8'hF8;
            16'd10056: data <= 8'h00;
            16'd10057: data <= 8'hF8;
            16'd10058: data <= 8'h00;
            16'd10059: data <= 8'hF8;
            16'd10060: data <= 8'h00;
            16'd10061: data <= 8'hF8;
            16'd10062: data <= 8'h00;
            16'd10063: data <= 8'hF8;
            16'd10064: data <= 8'h00;
            16'd10065: data <= 8'hF8;
            16'd10066: data <= 8'h00;
            16'd10067: data <= 8'hF8;
            16'd10068: data <= 8'h00;
            16'd10069: data <= 8'hF8;
            16'd10070: data <= 8'h00;
            16'd10071: data <= 8'hF8;
            16'd10072: data <= 8'h00;
            16'd10073: data <= 8'hF8;
            16'd10074: data <= 8'h00;
            16'd10075: data <= 8'hF8;
            16'd10076: data <= 8'h00;
            16'd10077: data <= 8'hF8;
            16'd10078: data <= 8'h00;
            16'd10079: data <= 8'hF8;
            16'd10080: data <= 8'hFF;
            16'd10081: data <= 8'hFF;
            16'd10082: data <= 8'h00;
            16'd10083: data <= 8'hF8;
            16'd10084: data <= 8'h00;
            16'd10085: data <= 8'hF8;
            16'd10086: data <= 8'h00;
            16'd10087: data <= 8'hF8;
            16'd10088: data <= 8'h00;
            16'd10089: data <= 8'hF8;
            16'd10090: data <= 8'h00;
            16'd10091: data <= 8'hF8;
            16'd10092: data <= 8'h00;
            16'd10093: data <= 8'hF8;
            16'd10094: data <= 8'h00;
            16'd10095: data <= 8'hF8;
            16'd10096: data <= 8'h00;
            16'd10097: data <= 8'hF8;
            16'd10098: data <= 8'h00;
            16'd10099: data <= 8'hF8;
            16'd10100: data <= 8'h00;
            16'd10101: data <= 8'hF8;
            16'd10102: data <= 8'h00;
            16'd10103: data <= 8'hF8;
            16'd10104: data <= 8'h00;
            16'd10105: data <= 8'hF8;
            16'd10106: data <= 8'h00;
            16'd10107: data <= 8'hF8;
            16'd10108: data <= 8'h00;
            16'd10109: data <= 8'hF8;
            16'd10110: data <= 8'h00;
            16'd10111: data <= 8'hF8;
            16'd10112: data <= 8'h00;
            16'd10113: data <= 8'hF8;
            16'd10114: data <= 8'h00;
            16'd10115: data <= 8'hF8;
            16'd10116: data <= 8'h00;
            16'd10117: data <= 8'hF8;
            16'd10118: data <= 8'h00;
            16'd10119: data <= 8'hF8;
            16'd10120: data <= 8'hFF;
            16'd10121: data <= 8'hFF;
            16'd10122: data <= 8'h00;
            16'd10123: data <= 8'hF8;
            16'd10124: data <= 8'h00;
            16'd10125: data <= 8'hF8;
            16'd10126: data <= 8'h00;
            16'd10127: data <= 8'hF8;
            16'd10128: data <= 8'h00;
            16'd10129: data <= 8'hF8;
            16'd10130: data <= 8'h00;
            16'd10131: data <= 8'hF8;
            16'd10132: data <= 8'h00;
            16'd10133: data <= 8'hF8;
            16'd10134: data <= 8'h00;
            16'd10135: data <= 8'hF8;
            16'd10136: data <= 8'h00;
            16'd10137: data <= 8'hF8;
            16'd10138: data <= 8'h00;
            16'd10139: data <= 8'hF8;
            16'd10140: data <= 8'h00;
            16'd10141: data <= 8'hF8;
            16'd10142: data <= 8'h00;
            16'd10143: data <= 8'hF8;
            16'd10144: data <= 8'h00;
            16'd10145: data <= 8'hF8;
            16'd10146: data <= 8'h00;
            16'd10147: data <= 8'hF8;
            16'd10148: data <= 8'h00;
            16'd10149: data <= 8'hF8;
            16'd10150: data <= 8'h00;
            16'd10151: data <= 8'hF8;
            16'd10152: data <= 8'h00;
            16'd10153: data <= 8'hF8;
            16'd10154: data <= 8'h00;
            16'd10155: data <= 8'hF8;
            16'd10156: data <= 8'h00;
            16'd10157: data <= 8'hF8;
            16'd10158: data <= 8'h00;
            16'd10159: data <= 8'hF8;
            16'd10160: data <= 8'hFF;
            16'd10161: data <= 8'hFF;
            16'd10162: data <= 8'h00;
            16'd10163: data <= 8'hF8;
            16'd10164: data <= 8'h00;
            16'd10165: data <= 8'hF8;
            16'd10166: data <= 8'h00;
            16'd10167: data <= 8'hF8;
            16'd10168: data <= 8'h00;
            16'd10169: data <= 8'hF8;
            16'd10170: data <= 8'h00;
            16'd10171: data <= 8'hF8;
            16'd10172: data <= 8'h00;
            16'd10173: data <= 8'hF8;
            16'd10174: data <= 8'h00;
            16'd10175: data <= 8'hF8;
            16'd10176: data <= 8'h00;
            16'd10177: data <= 8'hF8;
            16'd10178: data <= 8'h00;
            16'd10179: data <= 8'hF8;
            16'd10180: data <= 8'h00;
            16'd10181: data <= 8'hF8;
            16'd10182: data <= 8'h00;
            16'd10183: data <= 8'hF8;
            16'd10184: data <= 8'h00;
            16'd10185: data <= 8'hF8;
            16'd10186: data <= 8'h00;
            16'd10187: data <= 8'hF8;
            16'd10188: data <= 8'h00;
            16'd10189: data <= 8'hF8;
            16'd10190: data <= 8'h00;
            16'd10191: data <= 8'hF8;
            16'd10192: data <= 8'h00;
            16'd10193: data <= 8'hF8;
            16'd10194: data <= 8'h00;
            16'd10195: data <= 8'hF8;
            16'd10196: data <= 8'h00;
            16'd10197: data <= 8'hF8;
            16'd10198: data <= 8'h00;
            16'd10199: data <= 8'hF8;
            16'd10200: data <= 8'hFF;
            16'd10201: data <= 8'hFF;
            16'd10202: data <= 8'h00;
            16'd10203: data <= 8'hF8;
            16'd10204: data <= 8'h00;
            16'd10205: data <= 8'hF8;
            16'd10206: data <= 8'h00;
            16'd10207: data <= 8'hF8;
            16'd10208: data <= 8'h00;
            16'd10209: data <= 8'hF8;
            16'd10210: data <= 8'h00;
            16'd10211: data <= 8'hF8;
            16'd10212: data <= 8'h00;
            16'd10213: data <= 8'hF8;
            16'd10214: data <= 8'h00;
            16'd10215: data <= 8'hF8;
            16'd10216: data <= 8'h00;
            16'd10217: data <= 8'hF8;
            16'd10218: data <= 8'h00;
            16'd10219: data <= 8'hF8;
            16'd10220: data <= 8'h00;
            16'd10221: data <= 8'hF8;
            16'd10222: data <= 8'h00;
            16'd10223: data <= 8'hF8;
            16'd10224: data <= 8'h00;
            16'd10225: data <= 8'hF8;
            16'd10226: data <= 8'h00;
            16'd10227: data <= 8'hF8;
            16'd10228: data <= 8'h00;
            16'd10229: data <= 8'hF8;
            16'd10230: data <= 8'h00;
            16'd10231: data <= 8'hF8;
            16'd10232: data <= 8'h00;
            16'd10233: data <= 8'hF8;
            16'd10234: data <= 8'h00;
            16'd10235: data <= 8'hF8;
            16'd10236: data <= 8'h00;
            16'd10237: data <= 8'hF8;
            16'd10238: data <= 8'h00;
            16'd10239: data <= 8'hF8;
            16'd10240: data <= 8'hFF;
            16'd10241: data <= 8'hFF;
            16'd10242: data <= 8'h00;
            16'd10243: data <= 8'hF8;
            16'd10244: data <= 8'h00;
            16'd10245: data <= 8'hF8;
            16'd10246: data <= 8'h00;
            16'd10247: data <= 8'hF8;
            16'd10248: data <= 8'h00;
            16'd10249: data <= 8'hF8;
            16'd10250: data <= 8'h00;
            16'd10251: data <= 8'hF8;
            16'd10252: data <= 8'h00;
            16'd10253: data <= 8'hF8;
            16'd10254: data <= 8'h00;
            16'd10255: data <= 8'hF8;
            16'd10256: data <= 8'h00;
            16'd10257: data <= 8'hF8;
            16'd10258: data <= 8'h00;
            16'd10259: data <= 8'hF8;
            16'd10260: data <= 8'h00;
            16'd10261: data <= 8'hF8;
            16'd10262: data <= 8'h00;
            16'd10263: data <= 8'hF8;
            16'd10264: data <= 8'h00;
            16'd10265: data <= 8'hF8;
            16'd10266: data <= 8'h00;
            16'd10267: data <= 8'hF8;
            16'd10268: data <= 8'h00;
            16'd10269: data <= 8'hF8;
            16'd10270: data <= 8'h00;
            16'd10271: data <= 8'hF8;
            16'd10272: data <= 8'h00;
            16'd10273: data <= 8'hF8;
            16'd10274: data <= 8'h00;
            16'd10275: data <= 8'hF8;
            16'd10276: data <= 8'h00;
            16'd10277: data <= 8'hF8;
            16'd10278: data <= 8'h00;
            16'd10279: data <= 8'hF8;
            16'd10280: data <= 8'hFF;
            16'd10281: data <= 8'hFF;
            16'd10282: data <= 8'h00;
            16'd10283: data <= 8'hF8;
            16'd10284: data <= 8'h00;
            16'd10285: data <= 8'hF8;
            16'd10286: data <= 8'h00;
            16'd10287: data <= 8'hF8;
            16'd10288: data <= 8'h00;
            16'd10289: data <= 8'hF8;
            16'd10290: data <= 8'h00;
            16'd10291: data <= 8'hF8;
            16'd10292: data <= 8'h00;
            16'd10293: data <= 8'hF8;
            16'd10294: data <= 8'h00;
            16'd10295: data <= 8'hF8;
            16'd10296: data <= 8'h00;
            16'd10297: data <= 8'hF8;
            16'd10298: data <= 8'h00;
            16'd10299: data <= 8'hF8;
            16'd10300: data <= 8'h00;
            16'd10301: data <= 8'hF8;
            16'd10302: data <= 8'h00;
            16'd10303: data <= 8'hF8;
            16'd10304: data <= 8'h00;
            16'd10305: data <= 8'hF8;
            16'd10306: data <= 8'h00;
            16'd10307: data <= 8'hF8;
            16'd10308: data <= 8'h00;
            16'd10309: data <= 8'hF8;
            16'd10310: data <= 8'h00;
            16'd10311: data <= 8'hF8;
            16'd10312: data <= 8'h00;
            16'd10313: data <= 8'hF8;
            16'd10314: data <= 8'h00;
            16'd10315: data <= 8'hF8;
            16'd10316: data <= 8'h00;
            16'd10317: data <= 8'hF8;
            16'd10318: data <= 8'h00;
            16'd10319: data <= 8'hF8;
            16'd10320: data <= 8'hFF;
            16'd10321: data <= 8'hFF;
            16'd10322: data <= 8'h00;
            16'd10323: data <= 8'hF8;
            16'd10324: data <= 8'h00;
            16'd10325: data <= 8'hF8;
            16'd10326: data <= 8'h00;
            16'd10327: data <= 8'hF8;
            16'd10328: data <= 8'h00;
            16'd10329: data <= 8'hF8;
            16'd10330: data <= 8'h00;
            16'd10331: data <= 8'hF8;
            16'd10332: data <= 8'h00;
            16'd10333: data <= 8'hF8;
            16'd10334: data <= 8'h00;
            16'd10335: data <= 8'hF8;
            16'd10336: data <= 8'h00;
            16'd10337: data <= 8'hF8;
            16'd10338: data <= 8'h00;
            16'd10339: data <= 8'hF8;
            16'd10340: data <= 8'h00;
            16'd10341: data <= 8'hF8;
            16'd10342: data <= 8'h00;
            16'd10343: data <= 8'hF8;
            16'd10344: data <= 8'h00;
            16'd10345: data <= 8'hF8;
            16'd10346: data <= 8'h00;
            16'd10347: data <= 8'hF8;
            16'd10348: data <= 8'h00;
            16'd10349: data <= 8'hF8;
            16'd10350: data <= 8'h00;
            16'd10351: data <= 8'hF8;
            16'd10352: data <= 8'h00;
            16'd10353: data <= 8'hF8;
            16'd10354: data <= 8'h00;
            16'd10355: data <= 8'hF8;
            16'd10356: data <= 8'h00;
            16'd10357: data <= 8'hF8;
            16'd10358: data <= 8'h00;
            16'd10359: data <= 8'hF8;
            16'd10360: data <= 8'hFF;
            16'd10361: data <= 8'hFF;
            16'd10362: data <= 8'h00;
            16'd10363: data <= 8'hF8;
            16'd10364: data <= 8'h00;
            16'd10365: data <= 8'hF8;
            16'd10366: data <= 8'h00;
            16'd10367: data <= 8'hF8;
            16'd10368: data <= 8'h00;
            16'd10369: data <= 8'hF8;
            16'd10370: data <= 8'h00;
            16'd10371: data <= 8'hF8;
            16'd10372: data <= 8'h00;
            16'd10373: data <= 8'hF8;
            16'd10374: data <= 8'h00;
            16'd10375: data <= 8'hF8;
            16'd10376: data <= 8'h00;
            16'd10377: data <= 8'hF8;
            16'd10378: data <= 8'h00;
            16'd10379: data <= 8'hF8;
            16'd10380: data <= 8'h00;
            16'd10381: data <= 8'hF8;
            16'd10382: data <= 8'h00;
            16'd10383: data <= 8'hF8;
            16'd10384: data <= 8'h00;
            16'd10385: data <= 8'hF8;
            16'd10386: data <= 8'h00;
            16'd10387: data <= 8'hF8;
            16'd10388: data <= 8'h00;
            16'd10389: data <= 8'hF8;
            16'd10390: data <= 8'h00;
            16'd10391: data <= 8'hF8;
            16'd10392: data <= 8'h00;
            16'd10393: data <= 8'hF8;
            16'd10394: data <= 8'h00;
            16'd10395: data <= 8'hF8;
            16'd10396: data <= 8'h00;
            16'd10397: data <= 8'hF8;
            16'd10398: data <= 8'h00;
            16'd10399: data <= 8'hF8;
            16'd10400: data <= 8'hFF;
            16'd10401: data <= 8'hFF;
            16'd10402: data <= 8'h00;
            16'd10403: data <= 8'hF8;
            16'd10404: data <= 8'h00;
            16'd10405: data <= 8'hF8;
            16'd10406: data <= 8'h00;
            16'd10407: data <= 8'hF8;
            16'd10408: data <= 8'h00;
            16'd10409: data <= 8'hF8;
            16'd10410: data <= 8'h00;
            16'd10411: data <= 8'hF8;
            16'd10412: data <= 8'h00;
            16'd10413: data <= 8'hF8;
            16'd10414: data <= 8'h00;
            16'd10415: data <= 8'hF8;
            16'd10416: data <= 8'h00;
            16'd10417: data <= 8'hF8;
            16'd10418: data <= 8'h00;
            16'd10419: data <= 8'hF8;
            16'd10420: data <= 8'h00;
            16'd10421: data <= 8'hF8;
            16'd10422: data <= 8'h00;
            16'd10423: data <= 8'hF8;
            16'd10424: data <= 8'h00;
            16'd10425: data <= 8'hF8;
            16'd10426: data <= 8'h00;
            16'd10427: data <= 8'hF8;
            16'd10428: data <= 8'h00;
            16'd10429: data <= 8'hF8;
            16'd10430: data <= 8'h00;
            16'd10431: data <= 8'hF8;
            16'd10432: data <= 8'h00;
            16'd10433: data <= 8'hF8;
            16'd10434: data <= 8'h00;
            16'd10435: data <= 8'hF8;
            16'd10436: data <= 8'h00;
            16'd10437: data <= 8'hF8;
            16'd10438: data <= 8'h00;
            16'd10439: data <= 8'hF8;
            16'd10440: data <= 8'hFF;
            16'd10441: data <= 8'hFF;
            16'd10442: data <= 8'h00;
            16'd10443: data <= 8'hF8;
            16'd10444: data <= 8'h00;
            16'd10445: data <= 8'hF8;
            16'd10446: data <= 8'h00;
            16'd10447: data <= 8'hF8;
            16'd10448: data <= 8'h00;
            16'd10449: data <= 8'hF8;
            16'd10450: data <= 8'h00;
            16'd10451: data <= 8'hF8;
            16'd10452: data <= 8'h00;
            16'd10453: data <= 8'hF8;
            16'd10454: data <= 8'h00;
            16'd10455: data <= 8'hF8;
            16'd10456: data <= 8'h00;
            16'd10457: data <= 8'hF8;
            16'd10458: data <= 8'h00;
            16'd10459: data <= 8'hF8;
            16'd10460: data <= 8'h00;
            16'd10461: data <= 8'hF8;
            16'd10462: data <= 8'h00;
            16'd10463: data <= 8'hF8;
            16'd10464: data <= 8'h00;
            16'd10465: data <= 8'hF8;
            16'd10466: data <= 8'h00;
            16'd10467: data <= 8'hF8;
            16'd10468: data <= 8'h00;
            16'd10469: data <= 8'hF8;
            16'd10470: data <= 8'h00;
            16'd10471: data <= 8'hF8;
            16'd10472: data <= 8'h00;
            16'd10473: data <= 8'hF8;
            16'd10474: data <= 8'h00;
            16'd10475: data <= 8'hF8;
            16'd10476: data <= 8'h00;
            16'd10477: data <= 8'hF8;
            16'd10478: data <= 8'h00;
            16'd10479: data <= 8'hF8;
            16'd10480: data <= 8'hFF;
            16'd10481: data <= 8'hFF;
            16'd10482: data <= 8'h00;
            16'd10483: data <= 8'hF8;
            16'd10484: data <= 8'h00;
            16'd10485: data <= 8'hF8;
            16'd10486: data <= 8'h00;
            16'd10487: data <= 8'hF8;
            16'd10488: data <= 8'h00;
            16'd10489: data <= 8'hF8;
            16'd10490: data <= 8'h00;
            16'd10491: data <= 8'hF8;
            16'd10492: data <= 8'h00;
            16'd10493: data <= 8'hF8;
            16'd10494: data <= 8'h00;
            16'd10495: data <= 8'hF8;
            16'd10496: data <= 8'h00;
            16'd10497: data <= 8'hF8;
            16'd10498: data <= 8'h00;
            16'd10499: data <= 8'hF8;
            16'd10500: data <= 8'h00;
            16'd10501: data <= 8'hF8;
            16'd10502: data <= 8'h00;
            16'd10503: data <= 8'hF8;
            16'd10504: data <= 8'h00;
            16'd10505: data <= 8'hF8;
            16'd10506: data <= 8'h00;
            16'd10507: data <= 8'hF8;
            16'd10508: data <= 8'h00;
            16'd10509: data <= 8'hF8;
            16'd10510: data <= 8'h00;
            16'd10511: data <= 8'hF8;
            16'd10512: data <= 8'h00;
            16'd10513: data <= 8'hF8;
            16'd10514: data <= 8'h00;
            16'd10515: data <= 8'hF8;
            16'd10516: data <= 8'h00;
            16'd10517: data <= 8'hF8;
            16'd10518: data <= 8'h00;
            16'd10519: data <= 8'hF8;
            16'd10520: data <= 8'hFF;
            16'd10521: data <= 8'hFF;
            16'd10522: data <= 8'h00;
            16'd10523: data <= 8'hF8;
            16'd10524: data <= 8'h00;
            16'd10525: data <= 8'hF8;
            16'd10526: data <= 8'h00;
            16'd10527: data <= 8'hF8;
            16'd10528: data <= 8'h00;
            16'd10529: data <= 8'hF8;
            16'd10530: data <= 8'h00;
            16'd10531: data <= 8'hF8;
            16'd10532: data <= 8'h00;
            16'd10533: data <= 8'hF8;
            16'd10534: data <= 8'h00;
            16'd10535: data <= 8'hF8;
            16'd10536: data <= 8'h00;
            16'd10537: data <= 8'hF8;
            16'd10538: data <= 8'h00;
            16'd10539: data <= 8'hF8;
            16'd10540: data <= 8'h00;
            16'd10541: data <= 8'hF8;
            16'd10542: data <= 8'h00;
            16'd10543: data <= 8'hF8;
            16'd10544: data <= 8'h00;
            16'd10545: data <= 8'hF8;
            16'd10546: data <= 8'h00;
            16'd10547: data <= 8'hF8;
            16'd10548: data <= 8'h00;
            16'd10549: data <= 8'hF8;
            16'd10550: data <= 8'h00;
            16'd10551: data <= 8'hF8;
            16'd10552: data <= 8'h00;
            16'd10553: data <= 8'hF8;
            16'd10554: data <= 8'h00;
            16'd10555: data <= 8'hF8;
            16'd10556: data <= 8'h00;
            16'd10557: data <= 8'hF8;
            16'd10558: data <= 8'h00;
            16'd10559: data <= 8'hF8;
            16'd10560: data <= 8'hFF;
            16'd10561: data <= 8'hFF;
            16'd10562: data <= 8'h00;
            16'd10563: data <= 8'hF8;
            16'd10564: data <= 8'h00;
            16'd10565: data <= 8'hF8;
            16'd10566: data <= 8'h00;
            16'd10567: data <= 8'hF8;
            16'd10568: data <= 8'h00;
            16'd10569: data <= 8'hF8;
            16'd10570: data <= 8'h00;
            16'd10571: data <= 8'hF8;
            16'd10572: data <= 8'h00;
            16'd10573: data <= 8'hF8;
            16'd10574: data <= 8'h00;
            16'd10575: data <= 8'hF8;
            16'd10576: data <= 8'h00;
            16'd10577: data <= 8'hF8;
            16'd10578: data <= 8'h00;
            16'd10579: data <= 8'hF8;
            16'd10580: data <= 8'h00;
            16'd10581: data <= 8'hF8;
            16'd10582: data <= 8'h00;
            16'd10583: data <= 8'hF8;
            16'd10584: data <= 8'h00;
            16'd10585: data <= 8'hF8;
            16'd10586: data <= 8'h00;
            16'd10587: data <= 8'hF8;
            16'd10588: data <= 8'h00;
            16'd10589: data <= 8'hF8;
            16'd10590: data <= 8'h00;
            16'd10591: data <= 8'hF8;
            16'd10592: data <= 8'h00;
            16'd10593: data <= 8'hF8;
            16'd10594: data <= 8'h00;
            16'd10595: data <= 8'hF8;
            16'd10596: data <= 8'h00;
            16'd10597: data <= 8'hF8;
            16'd10598: data <= 8'h00;
            16'd10599: data <= 8'hF8;
            16'd10600: data <= 8'hFF;
            16'd10601: data <= 8'hFF;
            16'd10602: data <= 8'h00;
            16'd10603: data <= 8'hF8;
            16'd10604: data <= 8'h00;
            16'd10605: data <= 8'hF8;
            16'd10606: data <= 8'h00;
            16'd10607: data <= 8'hF8;
            16'd10608: data <= 8'h00;
            16'd10609: data <= 8'hF8;
            16'd10610: data <= 8'h00;
            16'd10611: data <= 8'hF8;
            16'd10612: data <= 8'h00;
            16'd10613: data <= 8'hF8;
            16'd10614: data <= 8'h00;
            16'd10615: data <= 8'hF8;
            16'd10616: data <= 8'h00;
            16'd10617: data <= 8'hF8;
            16'd10618: data <= 8'h00;
            16'd10619: data <= 8'hF8;
            16'd10620: data <= 8'h00;
            16'd10621: data <= 8'hF8;
            16'd10622: data <= 8'h00;
            16'd10623: data <= 8'hF8;
            16'd10624: data <= 8'h00;
            16'd10625: data <= 8'hF8;
            16'd10626: data <= 8'h00;
            16'd10627: data <= 8'hF8;
            16'd10628: data <= 8'h00;
            16'd10629: data <= 8'hF8;
            16'd10630: data <= 8'h00;
            16'd10631: data <= 8'hF8;
            16'd10632: data <= 8'h00;
            16'd10633: data <= 8'hF8;
            16'd10634: data <= 8'h00;
            16'd10635: data <= 8'hF8;
            16'd10636: data <= 8'h00;
            16'd10637: data <= 8'hF8;
            16'd10638: data <= 8'h00;
            16'd10639: data <= 8'hF8;
            16'd10640: data <= 8'hFF;
            16'd10641: data <= 8'hFF;
            16'd10642: data <= 8'h00;
            16'd10643: data <= 8'hF8;
            16'd10644: data <= 8'h00;
            16'd10645: data <= 8'hF8;
            16'd10646: data <= 8'h00;
            16'd10647: data <= 8'hF8;
            16'd10648: data <= 8'h00;
            16'd10649: data <= 8'hF8;
            16'd10650: data <= 8'h00;
            16'd10651: data <= 8'hF8;
            16'd10652: data <= 8'h00;
            16'd10653: data <= 8'hF8;
            16'd10654: data <= 8'h00;
            16'd10655: data <= 8'hF8;
            16'd10656: data <= 8'h00;
            16'd10657: data <= 8'hF8;
            16'd10658: data <= 8'h00;
            16'd10659: data <= 8'hF8;
            16'd10660: data <= 8'h00;
            16'd10661: data <= 8'hF8;
            16'd10662: data <= 8'h00;
            16'd10663: data <= 8'hF8;
            16'd10664: data <= 8'h00;
            16'd10665: data <= 8'hF8;
            16'd10666: data <= 8'h00;
            16'd10667: data <= 8'hF8;
            16'd10668: data <= 8'h00;
            16'd10669: data <= 8'hF8;
            16'd10670: data <= 8'h00;
            16'd10671: data <= 8'hF8;
            16'd10672: data <= 8'h00;
            16'd10673: data <= 8'hF8;
            16'd10674: data <= 8'h00;
            16'd10675: data <= 8'hF8;
            16'd10676: data <= 8'h00;
            16'd10677: data <= 8'hF8;
            16'd10678: data <= 8'h00;
            16'd10679: data <= 8'hF8;
            16'd10680: data <= 8'hFF;
            16'd10681: data <= 8'hFF;
            16'd10682: data <= 8'h00;
            16'd10683: data <= 8'hF8;
            16'd10684: data <= 8'h00;
            16'd10685: data <= 8'hF8;
            16'd10686: data <= 8'h00;
            16'd10687: data <= 8'hF8;
            16'd10688: data <= 8'h00;
            16'd10689: data <= 8'hF8;
            16'd10690: data <= 8'h00;
            16'd10691: data <= 8'hF8;
            16'd10692: data <= 8'h00;
            16'd10693: data <= 8'hF8;
            16'd10694: data <= 8'h00;
            16'd10695: data <= 8'hF8;
            16'd10696: data <= 8'h00;
            16'd10697: data <= 8'hF8;
            16'd10698: data <= 8'h00;
            16'd10699: data <= 8'hF8;
            16'd10700: data <= 8'h00;
            16'd10701: data <= 8'hF8;
            16'd10702: data <= 8'h00;
            16'd10703: data <= 8'hF8;
            16'd10704: data <= 8'h00;
            16'd10705: data <= 8'hF8;
            16'd10706: data <= 8'h00;
            16'd10707: data <= 8'hF8;
            16'd10708: data <= 8'h00;
            16'd10709: data <= 8'hF8;
            16'd10710: data <= 8'h00;
            16'd10711: data <= 8'hF8;
            16'd10712: data <= 8'h00;
            16'd10713: data <= 8'hF8;
            16'd10714: data <= 8'h00;
            16'd10715: data <= 8'hF8;
            16'd10716: data <= 8'h00;
            16'd10717: data <= 8'hF8;
            16'd10718: data <= 8'h00;
            16'd10719: data <= 8'hF8;
            16'd10720: data <= 8'hFF;
            16'd10721: data <= 8'hFF;
            16'd10722: data <= 8'h00;
            16'd10723: data <= 8'hF8;
            16'd10724: data <= 8'h00;
            16'd10725: data <= 8'hF8;
            16'd10726: data <= 8'h00;
            16'd10727: data <= 8'hF8;
            16'd10728: data <= 8'h00;
            16'd10729: data <= 8'hF8;
            16'd10730: data <= 8'h00;
            16'd10731: data <= 8'hF8;
            16'd10732: data <= 8'h00;
            16'd10733: data <= 8'hF8;
            16'd10734: data <= 8'h00;
            16'd10735: data <= 8'hF8;
            16'd10736: data <= 8'h00;
            16'd10737: data <= 8'hF8;
            16'd10738: data <= 8'h00;
            16'd10739: data <= 8'hF8;
            16'd10740: data <= 8'h00;
            16'd10741: data <= 8'hF8;
            16'd10742: data <= 8'h00;
            16'd10743: data <= 8'hF8;
            16'd10744: data <= 8'h00;
            16'd10745: data <= 8'hF8;
            16'd10746: data <= 8'h00;
            16'd10747: data <= 8'hF8;
            16'd10748: data <= 8'h00;
            16'd10749: data <= 8'hF8;
            16'd10750: data <= 8'h00;
            16'd10751: data <= 8'hF8;
            16'd10752: data <= 8'h00;
            16'd10753: data <= 8'hF8;
            16'd10754: data <= 8'h00;
            16'd10755: data <= 8'hF8;
            16'd10756: data <= 8'h00;
            16'd10757: data <= 8'hF8;
            16'd10758: data <= 8'h00;
            16'd10759: data <= 8'hF8;
            16'd10760: data <= 8'hFF;
            16'd10761: data <= 8'hFF;
            16'd10762: data <= 8'h00;
            16'd10763: data <= 8'hF8;
            16'd10764: data <= 8'h00;
            16'd10765: data <= 8'hF8;
            16'd10766: data <= 8'h00;
            16'd10767: data <= 8'hF8;
            16'd10768: data <= 8'h00;
            16'd10769: data <= 8'hF8;
            16'd10770: data <= 8'h00;
            16'd10771: data <= 8'hF8;
            16'd10772: data <= 8'h00;
            16'd10773: data <= 8'hF8;
            16'd10774: data <= 8'h00;
            16'd10775: data <= 8'hF8;
            16'd10776: data <= 8'h00;
            16'd10777: data <= 8'hF8;
            16'd10778: data <= 8'h00;
            16'd10779: data <= 8'hF8;
            16'd10780: data <= 8'h00;
            16'd10781: data <= 8'hF8;
            16'd10782: data <= 8'h00;
            16'd10783: data <= 8'hF8;
            16'd10784: data <= 8'h00;
            16'd10785: data <= 8'hF8;
            16'd10786: data <= 8'h00;
            16'd10787: data <= 8'hF8;
            16'd10788: data <= 8'h00;
            16'd10789: data <= 8'hF8;
            16'd10790: data <= 8'h00;
            16'd10791: data <= 8'hF8;
            16'd10792: data <= 8'h00;
            16'd10793: data <= 8'hF8;
            16'd10794: data <= 8'h00;
            16'd10795: data <= 8'hF8;
            16'd10796: data <= 8'h00;
            16'd10797: data <= 8'hF8;
            16'd10798: data <= 8'h00;
            16'd10799: data <= 8'hF8;
            16'd10800: data <= 8'hFF;
            16'd10801: data <= 8'hFF;
            16'd10802: data <= 8'h00;
            16'd10803: data <= 8'hF8;
            16'd10804: data <= 8'h00;
            16'd10805: data <= 8'hF8;
            16'd10806: data <= 8'h00;
            16'd10807: data <= 8'hF8;
            16'd10808: data <= 8'h00;
            16'd10809: data <= 8'hF8;
            16'd10810: data <= 8'h00;
            16'd10811: data <= 8'hF8;
            16'd10812: data <= 8'h00;
            16'd10813: data <= 8'hF8;
            16'd10814: data <= 8'h00;
            16'd10815: data <= 8'hF8;
            16'd10816: data <= 8'h00;
            16'd10817: data <= 8'hF8;
            16'd10818: data <= 8'h00;
            16'd10819: data <= 8'hF8;
            16'd10820: data <= 8'h00;
            16'd10821: data <= 8'hF8;
            16'd10822: data <= 8'h00;
            16'd10823: data <= 8'hF8;
            16'd10824: data <= 8'h00;
            16'd10825: data <= 8'hF8;
            16'd10826: data <= 8'h00;
            16'd10827: data <= 8'hF8;
            16'd10828: data <= 8'h00;
            16'd10829: data <= 8'hF8;
            16'd10830: data <= 8'h00;
            16'd10831: data <= 8'hF8;
            16'd10832: data <= 8'h00;
            16'd10833: data <= 8'hF8;
            16'd10834: data <= 8'h00;
            16'd10835: data <= 8'hF8;
            16'd10836: data <= 8'h00;
            16'd10837: data <= 8'hF8;
            16'd10838: data <= 8'h00;
            16'd10839: data <= 8'hF8;
            16'd10840: data <= 8'hFF;
            16'd10841: data <= 8'hFF;
            16'd10842: data <= 8'h00;
            16'd10843: data <= 8'hF8;
            16'd10844: data <= 8'h00;
            16'd10845: data <= 8'hF8;
            16'd10846: data <= 8'h00;
            16'd10847: data <= 8'hF8;
            16'd10848: data <= 8'h00;
            16'd10849: data <= 8'hF8;
            16'd10850: data <= 8'h00;
            16'd10851: data <= 8'hF8;
            16'd10852: data <= 8'h00;
            16'd10853: data <= 8'hF8;
            16'd10854: data <= 8'h00;
            16'd10855: data <= 8'hF8;
            16'd10856: data <= 8'h00;
            16'd10857: data <= 8'hF8;
            16'd10858: data <= 8'h00;
            16'd10859: data <= 8'hF8;
            16'd10860: data <= 8'h00;
            16'd10861: data <= 8'hF8;
            16'd10862: data <= 8'h00;
            16'd10863: data <= 8'hF8;
            16'd10864: data <= 8'h00;
            16'd10865: data <= 8'hF8;
            16'd10866: data <= 8'h00;
            16'd10867: data <= 8'hF8;
            16'd10868: data <= 8'h00;
            16'd10869: data <= 8'hF8;
            16'd10870: data <= 8'h00;
            16'd10871: data <= 8'hF8;
            16'd10872: data <= 8'h00;
            16'd10873: data <= 8'hF8;
            16'd10874: data <= 8'h00;
            16'd10875: data <= 8'hF8;
            16'd10876: data <= 8'h00;
            16'd10877: data <= 8'hF8;
            16'd10878: data <= 8'h00;
            16'd10879: data <= 8'hF8;
            16'd10880: data <= 8'hFF;
            16'd10881: data <= 8'hFF;
            16'd10882: data <= 8'h00;
            16'd10883: data <= 8'hF8;
            16'd10884: data <= 8'h00;
            16'd10885: data <= 8'hF8;
            16'd10886: data <= 8'h00;
            16'd10887: data <= 8'hF8;
            16'd10888: data <= 8'h00;
            16'd10889: data <= 8'hF8;
            16'd10890: data <= 8'h00;
            16'd10891: data <= 8'hF8;
            16'd10892: data <= 8'h00;
            16'd10893: data <= 8'hF8;
            16'd10894: data <= 8'h00;
            16'd10895: data <= 8'hF8;
            16'd10896: data <= 8'h00;
            16'd10897: data <= 8'hF8;
            16'd10898: data <= 8'h00;
            16'd10899: data <= 8'hF8;
            16'd10900: data <= 8'h00;
            16'd10901: data <= 8'hF8;
            16'd10902: data <= 8'h00;
            16'd10903: data <= 8'hF8;
            16'd10904: data <= 8'h00;
            16'd10905: data <= 8'hF8;
            16'd10906: data <= 8'h00;
            16'd10907: data <= 8'hF8;
            16'd10908: data <= 8'h00;
            16'd10909: data <= 8'hF8;
            16'd10910: data <= 8'h00;
            16'd10911: data <= 8'hF8;
            16'd10912: data <= 8'h00;
            16'd10913: data <= 8'hF8;
            16'd10914: data <= 8'h00;
            16'd10915: data <= 8'hF8;
            16'd10916: data <= 8'h00;
            16'd10917: data <= 8'hF8;
            16'd10918: data <= 8'h00;
            16'd10919: data <= 8'hF8;
            16'd10920: data <= 8'hFF;
            16'd10921: data <= 8'hFF;
            16'd10922: data <= 8'h00;
            16'd10923: data <= 8'hF8;
            16'd10924: data <= 8'h00;
            16'd10925: data <= 8'hF8;
            16'd10926: data <= 8'h00;
            16'd10927: data <= 8'hF8;
            16'd10928: data <= 8'h00;
            16'd10929: data <= 8'hF8;
            16'd10930: data <= 8'h00;
            16'd10931: data <= 8'hF8;
            16'd10932: data <= 8'h00;
            16'd10933: data <= 8'hF8;
            16'd10934: data <= 8'h00;
            16'd10935: data <= 8'hF8;
            16'd10936: data <= 8'h00;
            16'd10937: data <= 8'hF8;
            16'd10938: data <= 8'h00;
            16'd10939: data <= 8'hF8;
            16'd10940: data <= 8'h00;
            16'd10941: data <= 8'hF8;
            16'd10942: data <= 8'h00;
            16'd10943: data <= 8'hF8;
            16'd10944: data <= 8'h00;
            16'd10945: data <= 8'hF8;
            16'd10946: data <= 8'h00;
            16'd10947: data <= 8'hF8;
            16'd10948: data <= 8'h00;
            16'd10949: data <= 8'hF8;
            16'd10950: data <= 8'h00;
            16'd10951: data <= 8'hF8;
            16'd10952: data <= 8'h00;
            16'd10953: data <= 8'hF8;
            16'd10954: data <= 8'h00;
            16'd10955: data <= 8'hF8;
            16'd10956: data <= 8'h00;
            16'd10957: data <= 8'hF8;
            16'd10958: data <= 8'h00;
            16'd10959: data <= 8'hF8;
            16'd10960: data <= 8'hFF;
            16'd10961: data <= 8'hFF;
            16'd10962: data <= 8'h00;
            16'd10963: data <= 8'hF8;
            16'd10964: data <= 8'h00;
            16'd10965: data <= 8'hF8;
            16'd10966: data <= 8'h00;
            16'd10967: data <= 8'hF8;
            16'd10968: data <= 8'h00;
            16'd10969: data <= 8'hF8;
            16'd10970: data <= 8'h00;
            16'd10971: data <= 8'hF8;
            16'd10972: data <= 8'h00;
            16'd10973: data <= 8'hF8;
            16'd10974: data <= 8'h00;
            16'd10975: data <= 8'hF8;
            16'd10976: data <= 8'h00;
            16'd10977: data <= 8'hF8;
            16'd10978: data <= 8'h00;
            16'd10979: data <= 8'hF8;
            16'd10980: data <= 8'h00;
            16'd10981: data <= 8'hF8;
            16'd10982: data <= 8'h00;
            16'd10983: data <= 8'hF8;
            16'd10984: data <= 8'h00;
            16'd10985: data <= 8'hF8;
            16'd10986: data <= 8'h00;
            16'd10987: data <= 8'hF8;
            16'd10988: data <= 8'h00;
            16'd10989: data <= 8'hF8;
            16'd10990: data <= 8'h00;
            16'd10991: data <= 8'hF8;
            16'd10992: data <= 8'h00;
            16'd10993: data <= 8'hF8;
            16'd10994: data <= 8'h00;
            16'd10995: data <= 8'hF8;
            16'd10996: data <= 8'h00;
            16'd10997: data <= 8'hF8;
            16'd10998: data <= 8'h00;
            16'd10999: data <= 8'hF8;
            16'd11000: data <= 8'hFF;
            16'd11001: data <= 8'hFF;
            16'd11002: data <= 8'h00;
            16'd11003: data <= 8'hF8;
            16'd11004: data <= 8'h00;
            16'd11005: data <= 8'hF8;
            16'd11006: data <= 8'h00;
            16'd11007: data <= 8'hF8;
            16'd11008: data <= 8'h00;
            16'd11009: data <= 8'hF8;
            16'd11010: data <= 8'h00;
            16'd11011: data <= 8'hF8;
            16'd11012: data <= 8'h00;
            16'd11013: data <= 8'hF8;
            16'd11014: data <= 8'h00;
            16'd11015: data <= 8'hF8;
            16'd11016: data <= 8'h00;
            16'd11017: data <= 8'hF8;
            16'd11018: data <= 8'h00;
            16'd11019: data <= 8'hF8;
            16'd11020: data <= 8'h00;
            16'd11021: data <= 8'hF8;
            16'd11022: data <= 8'h00;
            16'd11023: data <= 8'hF8;
            16'd11024: data <= 8'h00;
            16'd11025: data <= 8'hF8;
            16'd11026: data <= 8'h00;
            16'd11027: data <= 8'hF8;
            16'd11028: data <= 8'h00;
            16'd11029: data <= 8'hF8;
            16'd11030: data <= 8'h00;
            16'd11031: data <= 8'hF8;
            16'd11032: data <= 8'h00;
            16'd11033: data <= 8'hF8;
            16'd11034: data <= 8'h00;
            16'd11035: data <= 8'hF8;
            16'd11036: data <= 8'h00;
            16'd11037: data <= 8'hF8;
            16'd11038: data <= 8'h00;
            16'd11039: data <= 8'hF8;
            16'd11040: data <= 8'hFF;
            16'd11041: data <= 8'hFF;
            16'd11042: data <= 8'h00;
            16'd11043: data <= 8'hF8;
            16'd11044: data <= 8'h00;
            16'd11045: data <= 8'hF8;
            16'd11046: data <= 8'h00;
            16'd11047: data <= 8'hF8;
            16'd11048: data <= 8'h00;
            16'd11049: data <= 8'hF8;
            16'd11050: data <= 8'h00;
            16'd11051: data <= 8'hF8;
            16'd11052: data <= 8'h00;
            16'd11053: data <= 8'hF8;
            16'd11054: data <= 8'h00;
            16'd11055: data <= 8'hF8;
            16'd11056: data <= 8'h00;
            16'd11057: data <= 8'hF8;
            16'd11058: data <= 8'h00;
            16'd11059: data <= 8'hF8;
            16'd11060: data <= 8'h00;
            16'd11061: data <= 8'hF8;
            16'd11062: data <= 8'h00;
            16'd11063: data <= 8'hF8;
            16'd11064: data <= 8'h00;
            16'd11065: data <= 8'hF8;
            16'd11066: data <= 8'h00;
            16'd11067: data <= 8'hF8;
            16'd11068: data <= 8'h00;
            16'd11069: data <= 8'hF8;
            16'd11070: data <= 8'h00;
            16'd11071: data <= 8'hF8;
            16'd11072: data <= 8'h00;
            16'd11073: data <= 8'hF8;
            16'd11074: data <= 8'h00;
            16'd11075: data <= 8'hF8;
            16'd11076: data <= 8'h00;
            16'd11077: data <= 8'hF8;
            16'd11078: data <= 8'h00;
            16'd11079: data <= 8'hF8;
            16'd11080: data <= 8'hFF;
            16'd11081: data <= 8'hFF;
            16'd11082: data <= 8'h00;
            16'd11083: data <= 8'hF8;
            16'd11084: data <= 8'h00;
            16'd11085: data <= 8'hF8;
            16'd11086: data <= 8'h00;
            16'd11087: data <= 8'hF8;
            16'd11088: data <= 8'h00;
            16'd11089: data <= 8'hF8;
            16'd11090: data <= 8'h00;
            16'd11091: data <= 8'hF8;
            16'd11092: data <= 8'h00;
            16'd11093: data <= 8'hF8;
            16'd11094: data <= 8'h00;
            16'd11095: data <= 8'hF8;
            16'd11096: data <= 8'h00;
            16'd11097: data <= 8'hF8;
            16'd11098: data <= 8'h00;
            16'd11099: data <= 8'hF8;
            16'd11100: data <= 8'h00;
            16'd11101: data <= 8'hF8;
            16'd11102: data <= 8'h00;
            16'd11103: data <= 8'hF8;
            16'd11104: data <= 8'h00;
            16'd11105: data <= 8'hF8;
            16'd11106: data <= 8'h00;
            16'd11107: data <= 8'hF8;
            16'd11108: data <= 8'h00;
            16'd11109: data <= 8'hF8;
            16'd11110: data <= 8'h00;
            16'd11111: data <= 8'hF8;
            16'd11112: data <= 8'h00;
            16'd11113: data <= 8'hF8;
            16'd11114: data <= 8'h00;
            16'd11115: data <= 8'hF8;
            16'd11116: data <= 8'h00;
            16'd11117: data <= 8'hF8;
            16'd11118: data <= 8'h00;
            16'd11119: data <= 8'hF8;
            16'd11120: data <= 8'hFF;
            16'd11121: data <= 8'hFF;
            16'd11122: data <= 8'h00;
            16'd11123: data <= 8'hF8;
            16'd11124: data <= 8'h00;
            16'd11125: data <= 8'hF8;
            16'd11126: data <= 8'h00;
            16'd11127: data <= 8'hF8;
            16'd11128: data <= 8'h00;
            16'd11129: data <= 8'hF8;
            16'd11130: data <= 8'h00;
            16'd11131: data <= 8'hF8;
            16'd11132: data <= 8'h00;
            16'd11133: data <= 8'hF8;
            16'd11134: data <= 8'h00;
            16'd11135: data <= 8'hF8;
            16'd11136: data <= 8'h00;
            16'd11137: data <= 8'hF8;
            16'd11138: data <= 8'h00;
            16'd11139: data <= 8'hF8;
            16'd11140: data <= 8'h00;
            16'd11141: data <= 8'hF8;
            16'd11142: data <= 8'h00;
            16'd11143: data <= 8'hF8;
            16'd11144: data <= 8'h00;
            16'd11145: data <= 8'hF8;
            16'd11146: data <= 8'h00;
            16'd11147: data <= 8'hF8;
            16'd11148: data <= 8'h00;
            16'd11149: data <= 8'hF8;
            16'd11150: data <= 8'h00;
            16'd11151: data <= 8'hF8;
            16'd11152: data <= 8'h00;
            16'd11153: data <= 8'hF8;
            16'd11154: data <= 8'h00;
            16'd11155: data <= 8'hF8;
            16'd11156: data <= 8'h00;
            16'd11157: data <= 8'hF8;
            16'd11158: data <= 8'h00;
            16'd11159: data <= 8'hF8;
            16'd11160: data <= 8'hFF;
            16'd11161: data <= 8'hFF;
            16'd11162: data <= 8'h00;
            16'd11163: data <= 8'hF8;
            16'd11164: data <= 8'h00;
            16'd11165: data <= 8'hF8;
            16'd11166: data <= 8'h00;
            16'd11167: data <= 8'hF8;
            16'd11168: data <= 8'h00;
            16'd11169: data <= 8'hF8;
            16'd11170: data <= 8'h00;
            16'd11171: data <= 8'hF8;
            16'd11172: data <= 8'h00;
            16'd11173: data <= 8'hF8;
            16'd11174: data <= 8'h00;
            16'd11175: data <= 8'hF8;
            16'd11176: data <= 8'h00;
            16'd11177: data <= 8'hF8;
            16'd11178: data <= 8'h00;
            16'd11179: data <= 8'hF8;
            16'd11180: data <= 8'h00;
            16'd11181: data <= 8'hF8;
            16'd11182: data <= 8'h00;
            16'd11183: data <= 8'hF8;
            16'd11184: data <= 8'h00;
            16'd11185: data <= 8'hF8;
            16'd11186: data <= 8'h00;
            16'd11187: data <= 8'hF8;
            16'd11188: data <= 8'h00;
            16'd11189: data <= 8'hF8;
            16'd11190: data <= 8'h00;
            16'd11191: data <= 8'hF8;
            16'd11192: data <= 8'h00;
            16'd11193: data <= 8'hF8;
            16'd11194: data <= 8'h00;
            16'd11195: data <= 8'hF8;
            16'd11196: data <= 8'h00;
            16'd11197: data <= 8'hF8;
            16'd11198: data <= 8'h00;
            16'd11199: data <= 8'hF8;
            16'd11200: data <= 8'hFF;
            16'd11201: data <= 8'hFF;
            16'd11202: data <= 8'h00;
            16'd11203: data <= 8'hF8;
            16'd11204: data <= 8'h00;
            16'd11205: data <= 8'hF8;
            16'd11206: data <= 8'h00;
            16'd11207: data <= 8'hF8;
            16'd11208: data <= 8'h00;
            16'd11209: data <= 8'hF8;
            16'd11210: data <= 8'h00;
            16'd11211: data <= 8'hF8;
            16'd11212: data <= 8'h00;
            16'd11213: data <= 8'hF8;
            16'd11214: data <= 8'h00;
            16'd11215: data <= 8'hF8;
            16'd11216: data <= 8'h00;
            16'd11217: data <= 8'hF8;
            16'd11218: data <= 8'h00;
            16'd11219: data <= 8'hF8;
            16'd11220: data <= 8'h00;
            16'd11221: data <= 8'hF8;
            16'd11222: data <= 8'h00;
            16'd11223: data <= 8'hF8;
            16'd11224: data <= 8'h00;
            16'd11225: data <= 8'hF8;
            16'd11226: data <= 8'h00;
            16'd11227: data <= 8'hF8;
            16'd11228: data <= 8'h00;
            16'd11229: data <= 8'hF8;
            16'd11230: data <= 8'h00;
            16'd11231: data <= 8'hF8;
            16'd11232: data <= 8'h00;
            16'd11233: data <= 8'hF8;
            16'd11234: data <= 8'h00;
            16'd11235: data <= 8'hF8;
            16'd11236: data <= 8'h00;
            16'd11237: data <= 8'hF8;
            16'd11238: data <= 8'h00;
            16'd11239: data <= 8'hF8;
            16'd11240: data <= 8'hFF;
            16'd11241: data <= 8'hFF;
            16'd11242: data <= 8'h00;
            16'd11243: data <= 8'hF8;
            16'd11244: data <= 8'h00;
            16'd11245: data <= 8'hF8;
            16'd11246: data <= 8'h00;
            16'd11247: data <= 8'hF8;
            16'd11248: data <= 8'h00;
            16'd11249: data <= 8'hF8;
            16'd11250: data <= 8'h00;
            16'd11251: data <= 8'hF8;
            16'd11252: data <= 8'h00;
            16'd11253: data <= 8'hF8;
            16'd11254: data <= 8'h00;
            16'd11255: data <= 8'hF8;
            16'd11256: data <= 8'h00;
            16'd11257: data <= 8'hF8;
            16'd11258: data <= 8'h00;
            16'd11259: data <= 8'hF8;
            16'd11260: data <= 8'h00;
            16'd11261: data <= 8'hF8;
            16'd11262: data <= 8'h00;
            16'd11263: data <= 8'hF8;
            16'd11264: data <= 8'h00;
            16'd11265: data <= 8'hF8;
            16'd11266: data <= 8'h00;
            16'd11267: data <= 8'hF8;
            16'd11268: data <= 8'h00;
            16'd11269: data <= 8'hF8;
            16'd11270: data <= 8'h00;
            16'd11271: data <= 8'hF8;
            16'd11272: data <= 8'h00;
            16'd11273: data <= 8'hF8;
            16'd11274: data <= 8'h00;
            16'd11275: data <= 8'hF8;
            16'd11276: data <= 8'h00;
            16'd11277: data <= 8'hF8;
            16'd11278: data <= 8'h00;
            16'd11279: data <= 8'hF8;
            16'd11280: data <= 8'hFF;
            16'd11281: data <= 8'hFF;
            16'd11282: data <= 8'h00;
            16'd11283: data <= 8'hF8;
            16'd11284: data <= 8'h00;
            16'd11285: data <= 8'hF8;
            16'd11286: data <= 8'h00;
            16'd11287: data <= 8'hF8;
            16'd11288: data <= 8'h00;
            16'd11289: data <= 8'hF8;
            16'd11290: data <= 8'h00;
            16'd11291: data <= 8'hF8;
            16'd11292: data <= 8'h00;
            16'd11293: data <= 8'hF8;
            16'd11294: data <= 8'h00;
            16'd11295: data <= 8'hF8;
            16'd11296: data <= 8'h00;
            16'd11297: data <= 8'hF8;
            16'd11298: data <= 8'h00;
            16'd11299: data <= 8'hF8;
            16'd11300: data <= 8'h00;
            16'd11301: data <= 8'hF8;
            16'd11302: data <= 8'h00;
            16'd11303: data <= 8'hF8;
            16'd11304: data <= 8'h00;
            16'd11305: data <= 8'hF8;
            16'd11306: data <= 8'h00;
            16'd11307: data <= 8'hF8;
            16'd11308: data <= 8'h00;
            16'd11309: data <= 8'hF8;
            16'd11310: data <= 8'h00;
            16'd11311: data <= 8'hF8;
            16'd11312: data <= 8'h00;
            16'd11313: data <= 8'hF8;
            16'd11314: data <= 8'h00;
            16'd11315: data <= 8'hF8;
            16'd11316: data <= 8'h00;
            16'd11317: data <= 8'hF8;
            16'd11318: data <= 8'h00;
            16'd11319: data <= 8'hF8;
            16'd11320: data <= 8'hFF;
            16'd11321: data <= 8'hFF;
            16'd11322: data <= 8'h00;
            16'd11323: data <= 8'hF8;
            16'd11324: data <= 8'h00;
            16'd11325: data <= 8'hF8;
            16'd11326: data <= 8'h00;
            16'd11327: data <= 8'hF8;
            16'd11328: data <= 8'h00;
            16'd11329: data <= 8'hF8;
            16'd11330: data <= 8'h00;
            16'd11331: data <= 8'hF8;
            16'd11332: data <= 8'h00;
            16'd11333: data <= 8'hF8;
            16'd11334: data <= 8'h00;
            16'd11335: data <= 8'hF8;
            16'd11336: data <= 8'h00;
            16'd11337: data <= 8'hF8;
            16'd11338: data <= 8'h00;
            16'd11339: data <= 8'hF8;
            16'd11340: data <= 8'h00;
            16'd11341: data <= 8'hF8;
            16'd11342: data <= 8'h00;
            16'd11343: data <= 8'hF8;
            16'd11344: data <= 8'h00;
            16'd11345: data <= 8'hF8;
            16'd11346: data <= 8'h00;
            16'd11347: data <= 8'hF8;
            16'd11348: data <= 8'h00;
            16'd11349: data <= 8'hF8;
            16'd11350: data <= 8'h00;
            16'd11351: data <= 8'hF8;
            16'd11352: data <= 8'h00;
            16'd11353: data <= 8'hF8;
            16'd11354: data <= 8'h00;
            16'd11355: data <= 8'hF8;
            16'd11356: data <= 8'h00;
            16'd11357: data <= 8'hF8;
            16'd11358: data <= 8'h00;
            16'd11359: data <= 8'hF8;
            16'd11360: data <= 8'hFF;
            16'd11361: data <= 8'hFF;
            16'd11362: data <= 8'h00;
            16'd11363: data <= 8'hF8;
            16'd11364: data <= 8'h00;
            16'd11365: data <= 8'hF8;
            16'd11366: data <= 8'h00;
            16'd11367: data <= 8'hF8;
            16'd11368: data <= 8'h00;
            16'd11369: data <= 8'hF8;
            16'd11370: data <= 8'h00;
            16'd11371: data <= 8'hF8;
            16'd11372: data <= 8'h00;
            16'd11373: data <= 8'hF8;
            16'd11374: data <= 8'h00;
            16'd11375: data <= 8'hF8;
            16'd11376: data <= 8'h00;
            16'd11377: data <= 8'hF8;
            16'd11378: data <= 8'h00;
            16'd11379: data <= 8'hF8;
            16'd11380: data <= 8'h00;
            16'd11381: data <= 8'hF8;
            16'd11382: data <= 8'h00;
            16'd11383: data <= 8'hF8;
            16'd11384: data <= 8'h00;
            16'd11385: data <= 8'hF8;
            16'd11386: data <= 8'h00;
            16'd11387: data <= 8'hF8;
            16'd11388: data <= 8'h00;
            16'd11389: data <= 8'hF8;
            16'd11390: data <= 8'h00;
            16'd11391: data <= 8'hF8;
            16'd11392: data <= 8'h00;
            16'd11393: data <= 8'hF8;
            16'd11394: data <= 8'h00;
            16'd11395: data <= 8'hF8;
            16'd11396: data <= 8'h00;
            16'd11397: data <= 8'hF8;
            16'd11398: data <= 8'h00;
            16'd11399: data <= 8'hF8;
            16'd11400: data <= 8'hFF;
            16'd11401: data <= 8'hFF;
            16'd11402: data <= 8'h00;
            16'd11403: data <= 8'hF8;
            16'd11404: data <= 8'h00;
            16'd11405: data <= 8'hF8;
            16'd11406: data <= 8'h00;
            16'd11407: data <= 8'hF8;
            16'd11408: data <= 8'h00;
            16'd11409: data <= 8'hF8;
            16'd11410: data <= 8'h00;
            16'd11411: data <= 8'hF8;
            16'd11412: data <= 8'h00;
            16'd11413: data <= 8'hF8;
            16'd11414: data <= 8'h00;
            16'd11415: data <= 8'hF8;
            16'd11416: data <= 8'h00;
            16'd11417: data <= 8'hF8;
            16'd11418: data <= 8'h00;
            16'd11419: data <= 8'hF8;
            16'd11420: data <= 8'h00;
            16'd11421: data <= 8'hF8;
            16'd11422: data <= 8'h00;
            16'd11423: data <= 8'hF8;
            16'd11424: data <= 8'h00;
            16'd11425: data <= 8'hF8;
            16'd11426: data <= 8'h00;
            16'd11427: data <= 8'hF8;
            16'd11428: data <= 8'h00;
            16'd11429: data <= 8'hF8;
            16'd11430: data <= 8'h00;
            16'd11431: data <= 8'hF8;
            16'd11432: data <= 8'h00;
            16'd11433: data <= 8'hF8;
            16'd11434: data <= 8'h00;
            16'd11435: data <= 8'hF8;
            16'd11436: data <= 8'h00;
            16'd11437: data <= 8'hF8;
            16'd11438: data <= 8'h00;
            16'd11439: data <= 8'hF8;
            16'd11440: data <= 8'hFF;
            16'd11441: data <= 8'hFF;
            16'd11442: data <= 8'h00;
            16'd11443: data <= 8'hF8;
            16'd11444: data <= 8'h00;
            16'd11445: data <= 8'hF8;
            16'd11446: data <= 8'h00;
            16'd11447: data <= 8'hF8;
            16'd11448: data <= 8'h00;
            16'd11449: data <= 8'hF8;
            16'd11450: data <= 8'h00;
            16'd11451: data <= 8'hF8;
            16'd11452: data <= 8'h00;
            16'd11453: data <= 8'hF8;
            16'd11454: data <= 8'h00;
            16'd11455: data <= 8'hF8;
            16'd11456: data <= 8'h00;
            16'd11457: data <= 8'hF8;
            16'd11458: data <= 8'h00;
            16'd11459: data <= 8'hF8;
            16'd11460: data <= 8'h00;
            16'd11461: data <= 8'hF8;
            16'd11462: data <= 8'h00;
            16'd11463: data <= 8'hF8;
            16'd11464: data <= 8'h00;
            16'd11465: data <= 8'hF8;
            16'd11466: data <= 8'h00;
            16'd11467: data <= 8'hF8;
            16'd11468: data <= 8'h00;
            16'd11469: data <= 8'hF8;
            16'd11470: data <= 8'h00;
            16'd11471: data <= 8'hF8;
            16'd11472: data <= 8'h00;
            16'd11473: data <= 8'hF8;
            16'd11474: data <= 8'h00;
            16'd11475: data <= 8'hF8;
            16'd11476: data <= 8'h00;
            16'd11477: data <= 8'hF8;
            16'd11478: data <= 8'h00;
            16'd11479: data <= 8'hF8;
            16'd11480: data <= 8'hFF;
            16'd11481: data <= 8'hFF;
            16'd11482: data <= 8'h00;
            16'd11483: data <= 8'hF8;
            16'd11484: data <= 8'h00;
            16'd11485: data <= 8'hF8;
            16'd11486: data <= 8'h00;
            16'd11487: data <= 8'hF8;
            16'd11488: data <= 8'h00;
            16'd11489: data <= 8'hF8;
            16'd11490: data <= 8'h00;
            16'd11491: data <= 8'hF8;
            16'd11492: data <= 8'h00;
            16'd11493: data <= 8'hF8;
            16'd11494: data <= 8'h00;
            16'd11495: data <= 8'hF8;
            16'd11496: data <= 8'h00;
            16'd11497: data <= 8'hF8;
            16'd11498: data <= 8'h00;
            16'd11499: data <= 8'hF8;
            16'd11500: data <= 8'h00;
            16'd11501: data <= 8'hF8;
            16'd11502: data <= 8'h00;
            16'd11503: data <= 8'hF8;
            16'd11504: data <= 8'h00;
            16'd11505: data <= 8'hF8;
            16'd11506: data <= 8'h00;
            16'd11507: data <= 8'hF8;
            16'd11508: data <= 8'h00;
            16'd11509: data <= 8'hF8;
            16'd11510: data <= 8'h00;
            16'd11511: data <= 8'hF8;
            16'd11512: data <= 8'h00;
            16'd11513: data <= 8'hF8;
            16'd11514: data <= 8'h00;
            16'd11515: data <= 8'hF8;
            16'd11516: data <= 8'h00;
            16'd11517: data <= 8'hF8;
            16'd11518: data <= 8'h00;
            16'd11519: data <= 8'hF8;
            16'd11520: data <= 8'hFF;
            16'd11521: data <= 8'hFF;
            16'd11522: data <= 8'h00;
            16'd11523: data <= 8'hF8;
            16'd11524: data <= 8'h00;
            16'd11525: data <= 8'hF8;
            16'd11526: data <= 8'h00;
            16'd11527: data <= 8'hF8;
            16'd11528: data <= 8'h00;
            16'd11529: data <= 8'hF8;
            16'd11530: data <= 8'h00;
            16'd11531: data <= 8'hF8;
            16'd11532: data <= 8'h00;
            16'd11533: data <= 8'hF8;
            16'd11534: data <= 8'h00;
            16'd11535: data <= 8'hF8;
            16'd11536: data <= 8'h00;
            16'd11537: data <= 8'hF8;
            16'd11538: data <= 8'h00;
            16'd11539: data <= 8'hF8;
            16'd11540: data <= 8'h00;
            16'd11541: data <= 8'hF8;
            16'd11542: data <= 8'h00;
            16'd11543: data <= 8'hF8;
            16'd11544: data <= 8'h00;
            16'd11545: data <= 8'hF8;
            16'd11546: data <= 8'h00;
            16'd11547: data <= 8'hF8;
            16'd11548: data <= 8'h00;
            16'd11549: data <= 8'hF8;
            16'd11550: data <= 8'h00;
            16'd11551: data <= 8'hF8;
            16'd11552: data <= 8'h00;
            16'd11553: data <= 8'hF8;
            16'd11554: data <= 8'h00;
            16'd11555: data <= 8'hF8;
            16'd11556: data <= 8'h00;
            16'd11557: data <= 8'hF8;
            16'd11558: data <= 8'h00;
            16'd11559: data <= 8'hF8;
            16'd11560: data <= 8'hFF;
            16'd11561: data <= 8'hFF;
            16'd11562: data <= 8'h00;
            16'd11563: data <= 8'hF8;
            16'd11564: data <= 8'h00;
            16'd11565: data <= 8'hF8;
            16'd11566: data <= 8'h00;
            16'd11567: data <= 8'hF8;
            16'd11568: data <= 8'h00;
            16'd11569: data <= 8'hF8;
            16'd11570: data <= 8'h00;
            16'd11571: data <= 8'hF8;
            16'd11572: data <= 8'h00;
            16'd11573: data <= 8'hF8;
            16'd11574: data <= 8'h00;
            16'd11575: data <= 8'hF8;
            16'd11576: data <= 8'h00;
            16'd11577: data <= 8'hF8;
            16'd11578: data <= 8'h00;
            16'd11579: data <= 8'hF8;
            16'd11580: data <= 8'h00;
            16'd11581: data <= 8'hF8;
            16'd11582: data <= 8'h00;
            16'd11583: data <= 8'hF8;
            16'd11584: data <= 8'h00;
            16'd11585: data <= 8'hF8;
            16'd11586: data <= 8'h00;
            16'd11587: data <= 8'hF8;
            16'd11588: data <= 8'h00;
            16'd11589: data <= 8'hF8;
            16'd11590: data <= 8'h00;
            16'd11591: data <= 8'hF8;
            16'd11592: data <= 8'h00;
            16'd11593: data <= 8'hF8;
            16'd11594: data <= 8'h00;
            16'd11595: data <= 8'hF8;
            16'd11596: data <= 8'h00;
            16'd11597: data <= 8'hF8;
            16'd11598: data <= 8'h00;
            16'd11599: data <= 8'hF8;
            16'd11600: data <= 8'hFF;
            16'd11601: data <= 8'hFF;
            16'd11602: data <= 8'h00;
            16'd11603: data <= 8'hF8;
            16'd11604: data <= 8'h00;
            16'd11605: data <= 8'hF8;
            16'd11606: data <= 8'h00;
            16'd11607: data <= 8'hF8;
            16'd11608: data <= 8'h00;
            16'd11609: data <= 8'hF8;
            16'd11610: data <= 8'h00;
            16'd11611: data <= 8'hF8;
            16'd11612: data <= 8'h00;
            16'd11613: data <= 8'hF8;
            16'd11614: data <= 8'h00;
            16'd11615: data <= 8'hF8;
            16'd11616: data <= 8'h00;
            16'd11617: data <= 8'hF8;
            16'd11618: data <= 8'h00;
            16'd11619: data <= 8'hF8;
            16'd11620: data <= 8'h00;
            16'd11621: data <= 8'hF8;
            16'd11622: data <= 8'h00;
            16'd11623: data <= 8'hF8;
            16'd11624: data <= 8'h00;
            16'd11625: data <= 8'hF8;
            16'd11626: data <= 8'h00;
            16'd11627: data <= 8'hF8;
            16'd11628: data <= 8'h00;
            16'd11629: data <= 8'hF8;
            16'd11630: data <= 8'h00;
            16'd11631: data <= 8'hF8;
            16'd11632: data <= 8'h00;
            16'd11633: data <= 8'hF8;
            16'd11634: data <= 8'h00;
            16'd11635: data <= 8'hF8;
            16'd11636: data <= 8'h00;
            16'd11637: data <= 8'hF8;
            16'd11638: data <= 8'h00;
            16'd11639: data <= 8'hF8;
            16'd11640: data <= 8'hFF;
            16'd11641: data <= 8'hFF;
            16'd11642: data <= 8'h00;
            16'd11643: data <= 8'hF8;
            16'd11644: data <= 8'h00;
            16'd11645: data <= 8'hF8;
            16'd11646: data <= 8'h00;
            16'd11647: data <= 8'hF8;
            16'd11648: data <= 8'h00;
            16'd11649: data <= 8'hF8;
            16'd11650: data <= 8'h00;
            16'd11651: data <= 8'hF8;
            16'd11652: data <= 8'h00;
            16'd11653: data <= 8'hF8;
            16'd11654: data <= 8'h00;
            16'd11655: data <= 8'hF8;
            16'd11656: data <= 8'h00;
            16'd11657: data <= 8'hF8;
            16'd11658: data <= 8'h00;
            16'd11659: data <= 8'hF8;
            16'd11660: data <= 8'h00;
            16'd11661: data <= 8'hF8;
            16'd11662: data <= 8'h00;
            16'd11663: data <= 8'hF8;
            16'd11664: data <= 8'h00;
            16'd11665: data <= 8'hF8;
            16'd11666: data <= 8'h00;
            16'd11667: data <= 8'hF8;
            16'd11668: data <= 8'h00;
            16'd11669: data <= 8'hF8;
            16'd11670: data <= 8'h00;
            16'd11671: data <= 8'hF8;
            16'd11672: data <= 8'h00;
            16'd11673: data <= 8'hF8;
            16'd11674: data <= 8'h00;
            16'd11675: data <= 8'hF8;
            16'd11676: data <= 8'h00;
            16'd11677: data <= 8'hF8;
            16'd11678: data <= 8'h00;
            16'd11679: data <= 8'hF8;
            16'd11680: data <= 8'hFF;
            16'd11681: data <= 8'hFF;
            16'd11682: data <= 8'h00;
            16'd11683: data <= 8'hF8;
            16'd11684: data <= 8'h00;
            16'd11685: data <= 8'hF8;
            16'd11686: data <= 8'h00;
            16'd11687: data <= 8'hF8;
            16'd11688: data <= 8'h00;
            16'd11689: data <= 8'hF8;
            16'd11690: data <= 8'h00;
            16'd11691: data <= 8'hF8;
            16'd11692: data <= 8'h00;
            16'd11693: data <= 8'hF8;
            16'd11694: data <= 8'h00;
            16'd11695: data <= 8'hF8;
            16'd11696: data <= 8'h00;
            16'd11697: data <= 8'hF8;
            16'd11698: data <= 8'h00;
            16'd11699: data <= 8'hF8;
            16'd11700: data <= 8'h00;
            16'd11701: data <= 8'hF8;
            16'd11702: data <= 8'h00;
            16'd11703: data <= 8'hF8;
            16'd11704: data <= 8'h00;
            16'd11705: data <= 8'hF8;
            16'd11706: data <= 8'h00;
            16'd11707: data <= 8'hF8;
            16'd11708: data <= 8'h00;
            16'd11709: data <= 8'hF8;
            16'd11710: data <= 8'h00;
            16'd11711: data <= 8'hF8;
            16'd11712: data <= 8'h00;
            16'd11713: data <= 8'hF8;
            16'd11714: data <= 8'h00;
            16'd11715: data <= 8'hF8;
            16'd11716: data <= 8'h00;
            16'd11717: data <= 8'hF8;
            16'd11718: data <= 8'h00;
            16'd11719: data <= 8'hF8;
            16'd11720: data <= 8'hFF;
            16'd11721: data <= 8'hFF;
            16'd11722: data <= 8'h00;
            16'd11723: data <= 8'hF8;
            16'd11724: data <= 8'h00;
            16'd11725: data <= 8'hF8;
            16'd11726: data <= 8'h00;
            16'd11727: data <= 8'hF8;
            16'd11728: data <= 8'h00;
            16'd11729: data <= 8'hF8;
            16'd11730: data <= 8'h00;
            16'd11731: data <= 8'hF8;
            16'd11732: data <= 8'h00;
            16'd11733: data <= 8'hF8;
            16'd11734: data <= 8'h00;
            16'd11735: data <= 8'hF8;
            16'd11736: data <= 8'h00;
            16'd11737: data <= 8'hF8;
            16'd11738: data <= 8'h00;
            16'd11739: data <= 8'hF8;
            16'd11740: data <= 8'h00;
            16'd11741: data <= 8'hF8;
            16'd11742: data <= 8'h00;
            16'd11743: data <= 8'hF8;
            16'd11744: data <= 8'h00;
            16'd11745: data <= 8'hF8;
            16'd11746: data <= 8'h00;
            16'd11747: data <= 8'hF8;
            16'd11748: data <= 8'h00;
            16'd11749: data <= 8'hF8;
            16'd11750: data <= 8'h00;
            16'd11751: data <= 8'hF8;
            16'd11752: data <= 8'h00;
            16'd11753: data <= 8'hF8;
            16'd11754: data <= 8'h00;
            16'd11755: data <= 8'hF8;
            16'd11756: data <= 8'h00;
            16'd11757: data <= 8'hF8;
            16'd11758: data <= 8'h00;
            16'd11759: data <= 8'hF8;
            16'd11760: data <= 8'hFF;
            16'd11761: data <= 8'hFF;
            16'd11762: data <= 8'h00;
            16'd11763: data <= 8'hF8;
            16'd11764: data <= 8'h00;
            16'd11765: data <= 8'hF8;
            16'd11766: data <= 8'h00;
            16'd11767: data <= 8'hF8;
            16'd11768: data <= 8'h00;
            16'd11769: data <= 8'hF8;
            16'd11770: data <= 8'h00;
            16'd11771: data <= 8'hF8;
            16'd11772: data <= 8'h00;
            16'd11773: data <= 8'hF8;
            16'd11774: data <= 8'h00;
            16'd11775: data <= 8'hF8;
            16'd11776: data <= 8'h00;
            16'd11777: data <= 8'hF8;
            16'd11778: data <= 8'h00;
            16'd11779: data <= 8'hF8;
            16'd11780: data <= 8'h00;
            16'd11781: data <= 8'hF8;
            16'd11782: data <= 8'h00;
            16'd11783: data <= 8'hF8;
            16'd11784: data <= 8'h00;
            16'd11785: data <= 8'hF8;
            16'd11786: data <= 8'h00;
            16'd11787: data <= 8'hF8;
            16'd11788: data <= 8'h00;
            16'd11789: data <= 8'hF8;
            16'd11790: data <= 8'h00;
            16'd11791: data <= 8'hF8;
            16'd11792: data <= 8'h00;
            16'd11793: data <= 8'hF8;
            16'd11794: data <= 8'h00;
            16'd11795: data <= 8'hF8;
            16'd11796: data <= 8'h00;
            16'd11797: data <= 8'hF8;
            16'd11798: data <= 8'h00;
            16'd11799: data <= 8'hF8;
            16'd11800: data <= 8'hFF;
            16'd11801: data <= 8'hFF;
            16'd11802: data <= 8'h00;
            16'd11803: data <= 8'hF8;
            16'd11804: data <= 8'h00;
            16'd11805: data <= 8'hF8;
            16'd11806: data <= 8'h00;
            16'd11807: data <= 8'hF8;
            16'd11808: data <= 8'h00;
            16'd11809: data <= 8'hF8;
            16'd11810: data <= 8'h00;
            16'd11811: data <= 8'hF8;
            16'd11812: data <= 8'h00;
            16'd11813: data <= 8'hF8;
            16'd11814: data <= 8'h00;
            16'd11815: data <= 8'hF8;
            16'd11816: data <= 8'h00;
            16'd11817: data <= 8'hF8;
            16'd11818: data <= 8'h00;
            16'd11819: data <= 8'hF8;
            16'd11820: data <= 8'h00;
            16'd11821: data <= 8'hF8;
            16'd11822: data <= 8'h00;
            16'd11823: data <= 8'hF8;
            16'd11824: data <= 8'h00;
            16'd11825: data <= 8'hF8;
            16'd11826: data <= 8'h00;
            16'd11827: data <= 8'hF8;
            16'd11828: data <= 8'h00;
            16'd11829: data <= 8'hF8;
            16'd11830: data <= 8'h00;
            16'd11831: data <= 8'hF8;
            16'd11832: data <= 8'h00;
            16'd11833: data <= 8'hF8;
            16'd11834: data <= 8'h00;
            16'd11835: data <= 8'hF8;
            16'd11836: data <= 8'h00;
            16'd11837: data <= 8'hF8;
            16'd11838: data <= 8'h00;
            16'd11839: data <= 8'hF8;
            16'd11840: data <= 8'hFF;
            16'd11841: data <= 8'hFF;
            16'd11842: data <= 8'h00;
            16'd11843: data <= 8'hF8;
            16'd11844: data <= 8'h00;
            16'd11845: data <= 8'hF8;
            16'd11846: data <= 8'h00;
            16'd11847: data <= 8'hF8;
            16'd11848: data <= 8'h00;
            16'd11849: data <= 8'hF8;
            16'd11850: data <= 8'h00;
            16'd11851: data <= 8'hF8;
            16'd11852: data <= 8'h00;
            16'd11853: data <= 8'hF8;
            16'd11854: data <= 8'h00;
            16'd11855: data <= 8'hF8;
            16'd11856: data <= 8'h00;
            16'd11857: data <= 8'hF8;
            16'd11858: data <= 8'h00;
            16'd11859: data <= 8'hF8;
            16'd11860: data <= 8'h00;
            16'd11861: data <= 8'hF8;
            16'd11862: data <= 8'h00;
            16'd11863: data <= 8'hF8;
            16'd11864: data <= 8'h00;
            16'd11865: data <= 8'hF8;
            16'd11866: data <= 8'h00;
            16'd11867: data <= 8'hF8;
            16'd11868: data <= 8'h00;
            16'd11869: data <= 8'hF8;
            16'd11870: data <= 8'h00;
            16'd11871: data <= 8'hF8;
            16'd11872: data <= 8'h00;
            16'd11873: data <= 8'hF8;
            16'd11874: data <= 8'h00;
            16'd11875: data <= 8'hF8;
            16'd11876: data <= 8'h00;
            16'd11877: data <= 8'hF8;
            16'd11878: data <= 8'h00;
            16'd11879: data <= 8'hF8;
            16'd11880: data <= 8'hFF;
            16'd11881: data <= 8'hFF;
            16'd11882: data <= 8'h00;
            16'd11883: data <= 8'hF8;
            16'd11884: data <= 8'h00;
            16'd11885: data <= 8'hF8;
            16'd11886: data <= 8'h00;
            16'd11887: data <= 8'hF8;
            16'd11888: data <= 8'h00;
            16'd11889: data <= 8'hF8;
            16'd11890: data <= 8'h00;
            16'd11891: data <= 8'hF8;
            16'd11892: data <= 8'h00;
            16'd11893: data <= 8'hF8;
            16'd11894: data <= 8'h00;
            16'd11895: data <= 8'hF8;
            16'd11896: data <= 8'h00;
            16'd11897: data <= 8'hF8;
            16'd11898: data <= 8'h00;
            16'd11899: data <= 8'hF8;
            16'd11900: data <= 8'h00;
            16'd11901: data <= 8'hF8;
            16'd11902: data <= 8'h00;
            16'd11903: data <= 8'hF8;
            16'd11904: data <= 8'h00;
            16'd11905: data <= 8'hF8;
            16'd11906: data <= 8'h00;
            16'd11907: data <= 8'hF8;
            16'd11908: data <= 8'h00;
            16'd11909: data <= 8'hF8;
            16'd11910: data <= 8'h00;
            16'd11911: data <= 8'hF8;
            16'd11912: data <= 8'h00;
            16'd11913: data <= 8'hF8;
            16'd11914: data <= 8'h00;
            16'd11915: data <= 8'hF8;
            16'd11916: data <= 8'h00;
            16'd11917: data <= 8'hF8;
            16'd11918: data <= 8'h00;
            16'd11919: data <= 8'hF8;
            16'd11920: data <= 8'hFF;
            16'd11921: data <= 8'hFF;
            16'd11922: data <= 8'h00;
            16'd11923: data <= 8'hF8;
            16'd11924: data <= 8'h00;
            16'd11925: data <= 8'hF8;
            16'd11926: data <= 8'h00;
            16'd11927: data <= 8'hF8;
            16'd11928: data <= 8'h00;
            16'd11929: data <= 8'hF8;
            16'd11930: data <= 8'h00;
            16'd11931: data <= 8'hF8;
            16'd11932: data <= 8'h00;
            16'd11933: data <= 8'hF8;
            16'd11934: data <= 8'h00;
            16'd11935: data <= 8'hF8;
            16'd11936: data <= 8'h00;
            16'd11937: data <= 8'hF8;
            16'd11938: data <= 8'h00;
            16'd11939: data <= 8'hF8;
            16'd11940: data <= 8'h00;
            16'd11941: data <= 8'hF8;
            16'd11942: data <= 8'h00;
            16'd11943: data <= 8'hF8;
            16'd11944: data <= 8'h00;
            16'd11945: data <= 8'hF8;
            16'd11946: data <= 8'h00;
            16'd11947: data <= 8'hF8;
            16'd11948: data <= 8'h00;
            16'd11949: data <= 8'hF8;
            16'd11950: data <= 8'h00;
            16'd11951: data <= 8'hF8;
            16'd11952: data <= 8'h00;
            16'd11953: data <= 8'hF8;
            16'd11954: data <= 8'h00;
            16'd11955: data <= 8'hF8;
            16'd11956: data <= 8'h00;
            16'd11957: data <= 8'hF8;
            16'd11958: data <= 8'h00;
            16'd11959: data <= 8'hF8;
            16'd11960: data <= 8'hFF;
            16'd11961: data <= 8'hFF;
            16'd11962: data <= 8'h00;
            16'd11963: data <= 8'hF8;
            16'd11964: data <= 8'h00;
            16'd11965: data <= 8'hF8;
            16'd11966: data <= 8'h00;
            16'd11967: data <= 8'hF8;
            16'd11968: data <= 8'h00;
            16'd11969: data <= 8'hF8;
            16'd11970: data <= 8'h00;
            16'd11971: data <= 8'hF8;
            16'd11972: data <= 8'h00;
            16'd11973: data <= 8'hF8;
            16'd11974: data <= 8'h00;
            16'd11975: data <= 8'hF8;
            16'd11976: data <= 8'h00;
            16'd11977: data <= 8'hF8;
            16'd11978: data <= 8'h00;
            16'd11979: data <= 8'hF8;
            16'd11980: data <= 8'h00;
            16'd11981: data <= 8'hF8;
            16'd11982: data <= 8'h00;
            16'd11983: data <= 8'hF8;
            16'd11984: data <= 8'h00;
            16'd11985: data <= 8'hF8;
            16'd11986: data <= 8'h00;
            16'd11987: data <= 8'hF8;
            16'd11988: data <= 8'h00;
            16'd11989: data <= 8'hF8;
            16'd11990: data <= 8'h00;
            16'd11991: data <= 8'hF8;
            16'd11992: data <= 8'h00;
            16'd11993: data <= 8'hF8;
            16'd11994: data <= 8'h00;
            16'd11995: data <= 8'hF8;
            16'd11996: data <= 8'h00;
            16'd11997: data <= 8'hF8;
            16'd11998: data <= 8'h00;
            16'd11999: data <= 8'hF8;
            16'd12000: data <= 8'hFF;
            16'd12001: data <= 8'hFF;
            16'd12002: data <= 8'h00;
            16'd12003: data <= 8'hF8;
            16'd12004: data <= 8'h00;
            16'd12005: data <= 8'hF8;
            16'd12006: data <= 8'h00;
            16'd12007: data <= 8'hF8;
            16'd12008: data <= 8'h00;
            16'd12009: data <= 8'hF8;
            16'd12010: data <= 8'h00;
            16'd12011: data <= 8'hF8;
            16'd12012: data <= 8'h00;
            16'd12013: data <= 8'hF8;
            16'd12014: data <= 8'h00;
            16'd12015: data <= 8'hF8;
            16'd12016: data <= 8'h00;
            16'd12017: data <= 8'hF8;
            16'd12018: data <= 8'h00;
            16'd12019: data <= 8'hF8;
            16'd12020: data <= 8'h00;
            16'd12021: data <= 8'hF8;
            16'd12022: data <= 8'h00;
            16'd12023: data <= 8'hF8;
            16'd12024: data <= 8'h00;
            16'd12025: data <= 8'hF8;
            16'd12026: data <= 8'h00;
            16'd12027: data <= 8'hF8;
            16'd12028: data <= 8'h00;
            16'd12029: data <= 8'hF8;
            16'd12030: data <= 8'h00;
            16'd12031: data <= 8'hF8;
            16'd12032: data <= 8'h00;
            16'd12033: data <= 8'hF8;
            16'd12034: data <= 8'h00;
            16'd12035: data <= 8'hF8;
            16'd12036: data <= 8'h00;
            16'd12037: data <= 8'hF8;
            16'd12038: data <= 8'h00;
            16'd12039: data <= 8'hF8;
            16'd12040: data <= 8'hFF;
            16'd12041: data <= 8'hFF;
            16'd12042: data <= 8'h00;
            16'd12043: data <= 8'hF8;
            16'd12044: data <= 8'h00;
            16'd12045: data <= 8'hF8;
            16'd12046: data <= 8'h00;
            16'd12047: data <= 8'hF8;
            16'd12048: data <= 8'h00;
            16'd12049: data <= 8'hF8;
            16'd12050: data <= 8'h00;
            16'd12051: data <= 8'hF8;
            16'd12052: data <= 8'h00;
            16'd12053: data <= 8'hF8;
            16'd12054: data <= 8'h00;
            16'd12055: data <= 8'hF8;
            16'd12056: data <= 8'h00;
            16'd12057: data <= 8'hF8;
            16'd12058: data <= 8'h00;
            16'd12059: data <= 8'hF8;
            16'd12060: data <= 8'h00;
            16'd12061: data <= 8'hF8;
            16'd12062: data <= 8'h00;
            16'd12063: data <= 8'hF8;
            16'd12064: data <= 8'h00;
            16'd12065: data <= 8'hF8;
            16'd12066: data <= 8'h00;
            16'd12067: data <= 8'hF8;
            16'd12068: data <= 8'h00;
            16'd12069: data <= 8'hF8;
            16'd12070: data <= 8'h00;
            16'd12071: data <= 8'hF8;
            16'd12072: data <= 8'h00;
            16'd12073: data <= 8'hF8;
            16'd12074: data <= 8'h00;
            16'd12075: data <= 8'hF8;
            16'd12076: data <= 8'h00;
            16'd12077: data <= 8'hF8;
            16'd12078: data <= 8'h00;
            16'd12079: data <= 8'hF8;
            16'd12080: data <= 8'hFF;
            16'd12081: data <= 8'hFF;
            16'd12082: data <= 8'h00;
            16'd12083: data <= 8'hF8;
            16'd12084: data <= 8'h00;
            16'd12085: data <= 8'hF8;
            16'd12086: data <= 8'h00;
            16'd12087: data <= 8'hF8;
            16'd12088: data <= 8'h00;
            16'd12089: data <= 8'hF8;
            16'd12090: data <= 8'h00;
            16'd12091: data <= 8'hF8;
            16'd12092: data <= 8'h00;
            16'd12093: data <= 8'hF8;
            16'd12094: data <= 8'h00;
            16'd12095: data <= 8'hF8;
            16'd12096: data <= 8'h00;
            16'd12097: data <= 8'hF8;
            16'd12098: data <= 8'h00;
            16'd12099: data <= 8'hF8;
            16'd12100: data <= 8'h00;
            16'd12101: data <= 8'hF8;
            16'd12102: data <= 8'h00;
            16'd12103: data <= 8'hF8;
            16'd12104: data <= 8'h00;
            16'd12105: data <= 8'hF8;
            16'd12106: data <= 8'h00;
            16'd12107: data <= 8'hF8;
            16'd12108: data <= 8'h00;
            16'd12109: data <= 8'hF8;
            16'd12110: data <= 8'h00;
            16'd12111: data <= 8'hF8;
            16'd12112: data <= 8'h00;
            16'd12113: data <= 8'hF8;
            16'd12114: data <= 8'h00;
            16'd12115: data <= 8'hF8;
            16'd12116: data <= 8'h00;
            16'd12117: data <= 8'hF8;
            16'd12118: data <= 8'h00;
            16'd12119: data <= 8'hF8;
            16'd12120: data <= 8'hFF;
            16'd12121: data <= 8'hFF;
            16'd12122: data <= 8'h00;
            16'd12123: data <= 8'hF8;
            16'd12124: data <= 8'h00;
            16'd12125: data <= 8'hF8;
            16'd12126: data <= 8'h00;
            16'd12127: data <= 8'hF8;
            16'd12128: data <= 8'h00;
            16'd12129: data <= 8'hF8;
            16'd12130: data <= 8'h00;
            16'd12131: data <= 8'hF8;
            16'd12132: data <= 8'h00;
            16'd12133: data <= 8'hF8;
            16'd12134: data <= 8'h00;
            16'd12135: data <= 8'hF8;
            16'd12136: data <= 8'h00;
            16'd12137: data <= 8'hF8;
            16'd12138: data <= 8'h00;
            16'd12139: data <= 8'hF8;
            16'd12140: data <= 8'h00;
            16'd12141: data <= 8'hF8;
            16'd12142: data <= 8'h00;
            16'd12143: data <= 8'hF8;
            16'd12144: data <= 8'h00;
            16'd12145: data <= 8'hF8;
            16'd12146: data <= 8'h00;
            16'd12147: data <= 8'hF8;
            16'd12148: data <= 8'h00;
            16'd12149: data <= 8'hF8;
            16'd12150: data <= 8'h00;
            16'd12151: data <= 8'hF8;
            16'd12152: data <= 8'h00;
            16'd12153: data <= 8'hF8;
            16'd12154: data <= 8'h00;
            16'd12155: data <= 8'hF8;
            16'd12156: data <= 8'h00;
            16'd12157: data <= 8'hF8;
            16'd12158: data <= 8'h00;
            16'd12159: data <= 8'hF8;
            16'd12160: data <= 8'hFF;
            16'd12161: data <= 8'hFF;
            16'd12162: data <= 8'h00;
            16'd12163: data <= 8'hF8;
            16'd12164: data <= 8'h00;
            16'd12165: data <= 8'hF8;
            16'd12166: data <= 8'h00;
            16'd12167: data <= 8'hF8;
            16'd12168: data <= 8'h00;
            16'd12169: data <= 8'hF8;
            16'd12170: data <= 8'h00;
            16'd12171: data <= 8'hF8;
            16'd12172: data <= 8'h00;
            16'd12173: data <= 8'hF8;
            16'd12174: data <= 8'h00;
            16'd12175: data <= 8'hF8;
            16'd12176: data <= 8'h00;
            16'd12177: data <= 8'hF8;
            16'd12178: data <= 8'h00;
            16'd12179: data <= 8'hF8;
            16'd12180: data <= 8'h00;
            16'd12181: data <= 8'hF8;
            16'd12182: data <= 8'h00;
            16'd12183: data <= 8'hF8;
            16'd12184: data <= 8'h00;
            16'd12185: data <= 8'hF8;
            16'd12186: data <= 8'h00;
            16'd12187: data <= 8'hF8;
            16'd12188: data <= 8'h00;
            16'd12189: data <= 8'hF8;
            16'd12190: data <= 8'h00;
            16'd12191: data <= 8'hF8;
            16'd12192: data <= 8'h00;
            16'd12193: data <= 8'hF8;
            16'd12194: data <= 8'h00;
            16'd12195: data <= 8'hF8;
            16'd12196: data <= 8'h00;
            16'd12197: data <= 8'hF8;
            16'd12198: data <= 8'h00;
            16'd12199: data <= 8'hF8;
            16'd12200: data <= 8'hFF;
            16'd12201: data <= 8'hFF;
            16'd12202: data <= 8'h00;
            16'd12203: data <= 8'hF8;
            16'd12204: data <= 8'h00;
            16'd12205: data <= 8'hF8;
            16'd12206: data <= 8'h00;
            16'd12207: data <= 8'hF8;
            16'd12208: data <= 8'h00;
            16'd12209: data <= 8'hF8;
            16'd12210: data <= 8'h00;
            16'd12211: data <= 8'hF8;
            16'd12212: data <= 8'h00;
            16'd12213: data <= 8'hF8;
            16'd12214: data <= 8'h00;
            16'd12215: data <= 8'hF8;
            16'd12216: data <= 8'h00;
            16'd12217: data <= 8'hF8;
            16'd12218: data <= 8'h00;
            16'd12219: data <= 8'hF8;
            16'd12220: data <= 8'h00;
            16'd12221: data <= 8'hF8;
            16'd12222: data <= 8'h00;
            16'd12223: data <= 8'hF8;
            16'd12224: data <= 8'h00;
            16'd12225: data <= 8'hF8;
            16'd12226: data <= 8'h00;
            16'd12227: data <= 8'hF8;
            16'd12228: data <= 8'h00;
            16'd12229: data <= 8'hF8;
            16'd12230: data <= 8'h00;
            16'd12231: data <= 8'hF8;
            16'd12232: data <= 8'h00;
            16'd12233: data <= 8'hF8;
            16'd12234: data <= 8'h00;
            16'd12235: data <= 8'hF8;
            16'd12236: data <= 8'h00;
            16'd12237: data <= 8'hF8;
            16'd12238: data <= 8'h00;
            16'd12239: data <= 8'hF8;
            16'd12240: data <= 8'hFF;
            16'd12241: data <= 8'hFF;
            16'd12242: data <= 8'h00;
            16'd12243: data <= 8'hF8;
            16'd12244: data <= 8'h00;
            16'd12245: data <= 8'hF8;
            16'd12246: data <= 8'h00;
            16'd12247: data <= 8'hF8;
            16'd12248: data <= 8'h00;
            16'd12249: data <= 8'hF8;
            16'd12250: data <= 8'h00;
            16'd12251: data <= 8'hF8;
            16'd12252: data <= 8'h00;
            16'd12253: data <= 8'hF8;
            16'd12254: data <= 8'h00;
            16'd12255: data <= 8'hF8;
            16'd12256: data <= 8'h00;
            16'd12257: data <= 8'hF8;
            16'd12258: data <= 8'h00;
            16'd12259: data <= 8'hF8;
            16'd12260: data <= 8'h00;
            16'd12261: data <= 8'hF8;
            16'd12262: data <= 8'h00;
            16'd12263: data <= 8'hF8;
            16'd12264: data <= 8'h00;
            16'd12265: data <= 8'hF8;
            16'd12266: data <= 8'h00;
            16'd12267: data <= 8'hF8;
            16'd12268: data <= 8'h00;
            16'd12269: data <= 8'hF8;
            16'd12270: data <= 8'h00;
            16'd12271: data <= 8'hF8;
            16'd12272: data <= 8'h00;
            16'd12273: data <= 8'hF8;
            16'd12274: data <= 8'h00;
            16'd12275: data <= 8'hF8;
            16'd12276: data <= 8'h00;
            16'd12277: data <= 8'hF8;
            16'd12278: data <= 8'h00;
            16'd12279: data <= 8'hF8;
            16'd12280: data <= 8'hFF;
            16'd12281: data <= 8'hFF;
            16'd12282: data <= 8'h00;
            16'd12283: data <= 8'hF8;
            16'd12284: data <= 8'h00;
            16'd12285: data <= 8'hF8;
            16'd12286: data <= 8'h00;
            16'd12287: data <= 8'hF8;
            16'd12288: data <= 8'h00;
            16'd12289: data <= 8'hF8;
            16'd12290: data <= 8'h00;
            16'd12291: data <= 8'hF8;
            16'd12292: data <= 8'h00;
            16'd12293: data <= 8'hF8;
            16'd12294: data <= 8'h00;
            16'd12295: data <= 8'hF8;
            16'd12296: data <= 8'h00;
            16'd12297: data <= 8'hF8;
            16'd12298: data <= 8'h00;
            16'd12299: data <= 8'hF8;
            16'd12300: data <= 8'h00;
            16'd12301: data <= 8'hF8;
            16'd12302: data <= 8'h00;
            16'd12303: data <= 8'hF8;
            16'd12304: data <= 8'h00;
            16'd12305: data <= 8'hF8;
            16'd12306: data <= 8'h00;
            16'd12307: data <= 8'hF8;
            16'd12308: data <= 8'h00;
            16'd12309: data <= 8'hF8;
            16'd12310: data <= 8'h00;
            16'd12311: data <= 8'hF8;
            16'd12312: data <= 8'h00;
            16'd12313: data <= 8'hF8;
            16'd12314: data <= 8'h00;
            16'd12315: data <= 8'hF8;
            16'd12316: data <= 8'h00;
            16'd12317: data <= 8'hF8;
            16'd12318: data <= 8'h00;
            16'd12319: data <= 8'hF8;
            16'd12320: data <= 8'hFF;
            16'd12321: data <= 8'hFF;
            16'd12322: data <= 8'h00;
            16'd12323: data <= 8'hF8;
            16'd12324: data <= 8'h00;
            16'd12325: data <= 8'hF8;
            16'd12326: data <= 8'h00;
            16'd12327: data <= 8'hF8;
            16'd12328: data <= 8'h00;
            16'd12329: data <= 8'hF8;
            16'd12330: data <= 8'h00;
            16'd12331: data <= 8'hF8;
            16'd12332: data <= 8'h00;
            16'd12333: data <= 8'hF8;
            16'd12334: data <= 8'h00;
            16'd12335: data <= 8'hF8;
            16'd12336: data <= 8'h00;
            16'd12337: data <= 8'hF8;
            16'd12338: data <= 8'h00;
            16'd12339: data <= 8'hF8;
            16'd12340: data <= 8'h00;
            16'd12341: data <= 8'hF8;
            16'd12342: data <= 8'h00;
            16'd12343: data <= 8'hF8;
            16'd12344: data <= 8'h00;
            16'd12345: data <= 8'hF8;
            16'd12346: data <= 8'h00;
            16'd12347: data <= 8'hF8;
            16'd12348: data <= 8'h00;
            16'd12349: data <= 8'hF8;
            16'd12350: data <= 8'h00;
            16'd12351: data <= 8'hF8;
            16'd12352: data <= 8'h00;
            16'd12353: data <= 8'hF8;
            16'd12354: data <= 8'h00;
            16'd12355: data <= 8'hF8;
            16'd12356: data <= 8'h00;
            16'd12357: data <= 8'hF8;
            16'd12358: data <= 8'h00;
            16'd12359: data <= 8'hF8;
            16'd12360: data <= 8'hFF;
            16'd12361: data <= 8'hFF;
            16'd12362: data <= 8'h00;
            16'd12363: data <= 8'hF8;
            16'd12364: data <= 8'h00;
            16'd12365: data <= 8'hF8;
            16'd12366: data <= 8'h00;
            16'd12367: data <= 8'hF8;
            16'd12368: data <= 8'h00;
            16'd12369: data <= 8'hF8;
            16'd12370: data <= 8'h00;
            16'd12371: data <= 8'hF8;
            16'd12372: data <= 8'h00;
            16'd12373: data <= 8'hF8;
            16'd12374: data <= 8'h00;
            16'd12375: data <= 8'hF8;
            16'd12376: data <= 8'h00;
            16'd12377: data <= 8'hF8;
            16'd12378: data <= 8'h00;
            16'd12379: data <= 8'hF8;
            16'd12380: data <= 8'h00;
            16'd12381: data <= 8'hF8;
            16'd12382: data <= 8'h00;
            16'd12383: data <= 8'hF8;
            16'd12384: data <= 8'h00;
            16'd12385: data <= 8'hF8;
            16'd12386: data <= 8'h00;
            16'd12387: data <= 8'hF8;
            16'd12388: data <= 8'h00;
            16'd12389: data <= 8'hF8;
            16'd12390: data <= 8'h00;
            16'd12391: data <= 8'hF8;
            16'd12392: data <= 8'h00;
            16'd12393: data <= 8'hF8;
            16'd12394: data <= 8'h00;
            16'd12395: data <= 8'hF8;
            16'd12396: data <= 8'h00;
            16'd12397: data <= 8'hF8;
            16'd12398: data <= 8'h00;
            16'd12399: data <= 8'hF8;
            16'd12400: data <= 8'hFF;
            16'd12401: data <= 8'hFF;
            16'd12402: data <= 8'h00;
            16'd12403: data <= 8'hF8;
            16'd12404: data <= 8'h00;
            16'd12405: data <= 8'hF8;
            16'd12406: data <= 8'h00;
            16'd12407: data <= 8'hF8;
            16'd12408: data <= 8'h00;
            16'd12409: data <= 8'hF8;
            16'd12410: data <= 8'h00;
            16'd12411: data <= 8'hF8;
            16'd12412: data <= 8'h00;
            16'd12413: data <= 8'hF8;
            16'd12414: data <= 8'h00;
            16'd12415: data <= 8'hF8;
            16'd12416: data <= 8'h00;
            16'd12417: data <= 8'hF8;
            16'd12418: data <= 8'h00;
            16'd12419: data <= 8'hF8;
            16'd12420: data <= 8'h00;
            16'd12421: data <= 8'hF8;
            16'd12422: data <= 8'h00;
            16'd12423: data <= 8'hF8;
            16'd12424: data <= 8'h00;
            16'd12425: data <= 8'hF8;
            16'd12426: data <= 8'h00;
            16'd12427: data <= 8'hF8;
            16'd12428: data <= 8'h00;
            16'd12429: data <= 8'hF8;
            16'd12430: data <= 8'h00;
            16'd12431: data <= 8'hF8;
            16'd12432: data <= 8'h00;
            16'd12433: data <= 8'hF8;
            16'd12434: data <= 8'h00;
            16'd12435: data <= 8'hF8;
            16'd12436: data <= 8'h00;
            16'd12437: data <= 8'hF8;
            16'd12438: data <= 8'h00;
            16'd12439: data <= 8'hF8;
            16'd12440: data <= 8'hFF;
            16'd12441: data <= 8'hFF;
            16'd12442: data <= 8'h00;
            16'd12443: data <= 8'hF8;
            16'd12444: data <= 8'h00;
            16'd12445: data <= 8'hF8;
            16'd12446: data <= 8'h00;
            16'd12447: data <= 8'hF8;
            16'd12448: data <= 8'h00;
            16'd12449: data <= 8'hF8;
            16'd12450: data <= 8'h00;
            16'd12451: data <= 8'hF8;
            16'd12452: data <= 8'h00;
            16'd12453: data <= 8'hF8;
            16'd12454: data <= 8'h00;
            16'd12455: data <= 8'hF8;
            16'd12456: data <= 8'h00;
            16'd12457: data <= 8'hF8;
            16'd12458: data <= 8'h00;
            16'd12459: data <= 8'hF8;
            16'd12460: data <= 8'h00;
            16'd12461: data <= 8'hF8;
            16'd12462: data <= 8'h00;
            16'd12463: data <= 8'hF8;
            16'd12464: data <= 8'h00;
            16'd12465: data <= 8'hF8;
            16'd12466: data <= 8'h00;
            16'd12467: data <= 8'hF8;
            16'd12468: data <= 8'h00;
            16'd12469: data <= 8'hF8;
            16'd12470: data <= 8'h00;
            16'd12471: data <= 8'hF8;
            16'd12472: data <= 8'h00;
            16'd12473: data <= 8'hF8;
            16'd12474: data <= 8'h00;
            16'd12475: data <= 8'hF8;
            16'd12476: data <= 8'h00;
            16'd12477: data <= 8'hF8;
            16'd12478: data <= 8'h00;
            16'd12479: data <= 8'hF8;
            16'd12480: data <= 8'hFF;
            16'd12481: data <= 8'hFF;
            16'd12482: data <= 8'h00;
            16'd12483: data <= 8'hF8;
            16'd12484: data <= 8'h00;
            16'd12485: data <= 8'hF8;
            16'd12486: data <= 8'h00;
            16'd12487: data <= 8'hF8;
            16'd12488: data <= 8'h00;
            16'd12489: data <= 8'hF8;
            16'd12490: data <= 8'h00;
            16'd12491: data <= 8'hF8;
            16'd12492: data <= 8'h00;
            16'd12493: data <= 8'hF8;
            16'd12494: data <= 8'h00;
            16'd12495: data <= 8'hF8;
            16'd12496: data <= 8'h00;
            16'd12497: data <= 8'hF8;
            16'd12498: data <= 8'h00;
            16'd12499: data <= 8'hF8;
            16'd12500: data <= 8'h00;
            16'd12501: data <= 8'hF8;
            16'd12502: data <= 8'h00;
            16'd12503: data <= 8'hF8;
            16'd12504: data <= 8'h00;
            16'd12505: data <= 8'hF8;
            16'd12506: data <= 8'h00;
            16'd12507: data <= 8'hF8;
            16'd12508: data <= 8'h00;
            16'd12509: data <= 8'hF8;
            16'd12510: data <= 8'h00;
            16'd12511: data <= 8'hF8;
            16'd12512: data <= 8'h00;
            16'd12513: data <= 8'hF8;
            16'd12514: data <= 8'h00;
            16'd12515: data <= 8'hF8;
            16'd12516: data <= 8'h00;
            16'd12517: data <= 8'hF8;
            16'd12518: data <= 8'h00;
            16'd12519: data <= 8'hF8;
            16'd12520: data <= 8'hFF;
            16'd12521: data <= 8'hFF;
            16'd12522: data <= 8'h00;
            16'd12523: data <= 8'hF8;
            16'd12524: data <= 8'h00;
            16'd12525: data <= 8'hF8;
            16'd12526: data <= 8'h00;
            16'd12527: data <= 8'hF8;
            16'd12528: data <= 8'h00;
            16'd12529: data <= 8'hF8;
            16'd12530: data <= 8'h00;
            16'd12531: data <= 8'hF8;
            16'd12532: data <= 8'h00;
            16'd12533: data <= 8'hF8;
            16'd12534: data <= 8'h00;
            16'd12535: data <= 8'hF8;
            16'd12536: data <= 8'h00;
            16'd12537: data <= 8'hF8;
            16'd12538: data <= 8'h00;
            16'd12539: data <= 8'hF8;
            16'd12540: data <= 8'h00;
            16'd12541: data <= 8'hF8;
            16'd12542: data <= 8'h00;
            16'd12543: data <= 8'hF8;
            16'd12544: data <= 8'h00;
            16'd12545: data <= 8'hF8;
            16'd12546: data <= 8'h00;
            16'd12547: data <= 8'hF8;
            16'd12548: data <= 8'h00;
            16'd12549: data <= 8'hF8;
            16'd12550: data <= 8'h00;
            16'd12551: data <= 8'hF8;
            16'd12552: data <= 8'h00;
            16'd12553: data <= 8'hF8;
            16'd12554: data <= 8'h00;
            16'd12555: data <= 8'hF8;
            16'd12556: data <= 8'h00;
            16'd12557: data <= 8'hF8;
            16'd12558: data <= 8'h00;
            16'd12559: data <= 8'hF8;
            16'd12560: data <= 8'hFF;
            16'd12561: data <= 8'hFF;
            16'd12562: data <= 8'h00;
            16'd12563: data <= 8'hF8;
            16'd12564: data <= 8'h00;
            16'd12565: data <= 8'hF8;
            16'd12566: data <= 8'h00;
            16'd12567: data <= 8'hF8;
            16'd12568: data <= 8'h00;
            16'd12569: data <= 8'hF8;
            16'd12570: data <= 8'h00;
            16'd12571: data <= 8'hF8;
            16'd12572: data <= 8'h00;
            16'd12573: data <= 8'hF8;
            16'd12574: data <= 8'h00;
            16'd12575: data <= 8'hF8;
            16'd12576: data <= 8'h00;
            16'd12577: data <= 8'hF8;
            16'd12578: data <= 8'h00;
            16'd12579: data <= 8'hF8;
            16'd12580: data <= 8'h00;
            16'd12581: data <= 8'hF8;
            16'd12582: data <= 8'h00;
            16'd12583: data <= 8'hF8;
            16'd12584: data <= 8'h00;
            16'd12585: data <= 8'hF8;
            16'd12586: data <= 8'h00;
            16'd12587: data <= 8'hF8;
            16'd12588: data <= 8'h00;
            16'd12589: data <= 8'hF8;
            16'd12590: data <= 8'h00;
            16'd12591: data <= 8'hF8;
            16'd12592: data <= 8'h00;
            16'd12593: data <= 8'hF8;
            16'd12594: data <= 8'h00;
            16'd12595: data <= 8'hF8;
            16'd12596: data <= 8'h00;
            16'd12597: data <= 8'hF8;
            16'd12598: data <= 8'h00;
            16'd12599: data <= 8'hF8;
            16'd12600: data <= 8'hFF;
            16'd12601: data <= 8'hFF;
            16'd12602: data <= 8'h00;
            16'd12603: data <= 8'hF8;
            16'd12604: data <= 8'h00;
            16'd12605: data <= 8'hF8;
            16'd12606: data <= 8'h00;
            16'd12607: data <= 8'hF8;
            16'd12608: data <= 8'h00;
            16'd12609: data <= 8'hF8;
            16'd12610: data <= 8'h00;
            16'd12611: data <= 8'hF8;
            16'd12612: data <= 8'h00;
            16'd12613: data <= 8'hF8;
            16'd12614: data <= 8'h00;
            16'd12615: data <= 8'hF8;
            16'd12616: data <= 8'h00;
            16'd12617: data <= 8'hF8;
            16'd12618: data <= 8'h00;
            16'd12619: data <= 8'hF8;
            16'd12620: data <= 8'h00;
            16'd12621: data <= 8'hF8;
            16'd12622: data <= 8'h00;
            16'd12623: data <= 8'hF8;
            16'd12624: data <= 8'h00;
            16'd12625: data <= 8'hF8;
            16'd12626: data <= 8'h00;
            16'd12627: data <= 8'hF8;
            16'd12628: data <= 8'h00;
            16'd12629: data <= 8'hF8;
            16'd12630: data <= 8'h00;
            16'd12631: data <= 8'hF8;
            16'd12632: data <= 8'h00;
            16'd12633: data <= 8'hF8;
            16'd12634: data <= 8'h00;
            16'd12635: data <= 8'hF8;
            16'd12636: data <= 8'h00;
            16'd12637: data <= 8'hF8;
            16'd12638: data <= 8'h00;
            16'd12639: data <= 8'hF8;
            16'd12640: data <= 8'hFF;
            16'd12641: data <= 8'hFF;
            16'd12642: data <= 8'h00;
            16'd12643: data <= 8'hF8;
            16'd12644: data <= 8'h00;
            16'd12645: data <= 8'hF8;
            16'd12646: data <= 8'h00;
            16'd12647: data <= 8'hF8;
            16'd12648: data <= 8'h00;
            16'd12649: data <= 8'hF8;
            16'd12650: data <= 8'h00;
            16'd12651: data <= 8'hF8;
            16'd12652: data <= 8'h00;
            16'd12653: data <= 8'hF8;
            16'd12654: data <= 8'h00;
            16'd12655: data <= 8'hF8;
            16'd12656: data <= 8'h00;
            16'd12657: data <= 8'hF8;
            16'd12658: data <= 8'h00;
            16'd12659: data <= 8'hF8;
            16'd12660: data <= 8'h00;
            16'd12661: data <= 8'hF8;
            16'd12662: data <= 8'h00;
            16'd12663: data <= 8'hF8;
            16'd12664: data <= 8'h00;
            16'd12665: data <= 8'hF8;
            16'd12666: data <= 8'h00;
            16'd12667: data <= 8'hF8;
            16'd12668: data <= 8'h00;
            16'd12669: data <= 8'hF8;
            16'd12670: data <= 8'h00;
            16'd12671: data <= 8'hF8;
            16'd12672: data <= 8'h00;
            16'd12673: data <= 8'hF8;
            16'd12674: data <= 8'h00;
            16'd12675: data <= 8'hF8;
            16'd12676: data <= 8'h00;
            16'd12677: data <= 8'hF8;
            16'd12678: data <= 8'h00;
            16'd12679: data <= 8'hF8;
            16'd12680: data <= 8'hFF;
            16'd12681: data <= 8'hFF;
            16'd12682: data <= 8'h00;
            16'd12683: data <= 8'hF8;
            16'd12684: data <= 8'h00;
            16'd12685: data <= 8'hF8;
            16'd12686: data <= 8'h00;
            16'd12687: data <= 8'hF8;
            16'd12688: data <= 8'h00;
            16'd12689: data <= 8'hF8;
            16'd12690: data <= 8'h00;
            16'd12691: data <= 8'hF8;
            16'd12692: data <= 8'h00;
            16'd12693: data <= 8'hF8;
            16'd12694: data <= 8'h00;
            16'd12695: data <= 8'hF8;
            16'd12696: data <= 8'h00;
            16'd12697: data <= 8'hF8;
            16'd12698: data <= 8'h00;
            16'd12699: data <= 8'hF8;
            16'd12700: data <= 8'h00;
            16'd12701: data <= 8'hF8;
            16'd12702: data <= 8'h00;
            16'd12703: data <= 8'hF8;
            16'd12704: data <= 8'h00;
            16'd12705: data <= 8'hF8;
            16'd12706: data <= 8'h00;
            16'd12707: data <= 8'hF8;
            16'd12708: data <= 8'h00;
            16'd12709: data <= 8'hF8;
            16'd12710: data <= 8'h00;
            16'd12711: data <= 8'hF8;
            16'd12712: data <= 8'h00;
            16'd12713: data <= 8'hF8;
            16'd12714: data <= 8'h00;
            16'd12715: data <= 8'hF8;
            16'd12716: data <= 8'h00;
            16'd12717: data <= 8'hF8;
            16'd12718: data <= 8'h00;
            16'd12719: data <= 8'hF8;
            16'd12720: data <= 8'hFF;
            16'd12721: data <= 8'hFF;
            16'd12722: data <= 8'hE0;
            16'd12723: data <= 8'h07;
            16'd12724: data <= 8'hE0;
            16'd12725: data <= 8'h07;
            16'd12726: data <= 8'hE0;
            16'd12727: data <= 8'h07;
            16'd12728: data <= 8'hE0;
            16'd12729: data <= 8'h07;
            16'd12730: data <= 8'hE0;
            16'd12731: data <= 8'h07;
            16'd12732: data <= 8'hE0;
            16'd12733: data <= 8'h07;
            16'd12734: data <= 8'hE0;
            16'd12735: data <= 8'h07;
            16'd12736: data <= 8'hE0;
            16'd12737: data <= 8'h07;
            16'd12738: data <= 8'hE0;
            16'd12739: data <= 8'h07;
            16'd12740: data <= 8'hE0;
            16'd12741: data <= 8'h07;
            16'd12742: data <= 8'hE0;
            16'd12743: data <= 8'h07;
            16'd12744: data <= 8'hE0;
            16'd12745: data <= 8'h07;
            16'd12746: data <= 8'hE0;
            16'd12747: data <= 8'h07;
            16'd12748: data <= 8'hE0;
            16'd12749: data <= 8'h07;
            16'd12750: data <= 8'hE0;
            16'd12751: data <= 8'h07;
            16'd12752: data <= 8'hE0;
            16'd12753: data <= 8'h07;
            16'd12754: data <= 8'hE0;
            16'd12755: data <= 8'h07;
            16'd12756: data <= 8'hE0;
            16'd12757: data <= 8'h07;
            16'd12758: data <= 8'hE0;
            16'd12759: data <= 8'h07;
            16'd12760: data <= 8'hFF;
            16'd12761: data <= 8'hFF;
            16'd12762: data <= 8'hE0;
            16'd12763: data <= 8'h07;
            16'd12764: data <= 8'hE0;
            16'd12765: data <= 8'h07;
            16'd12766: data <= 8'hE0;
            16'd12767: data <= 8'h07;
            16'd12768: data <= 8'hE0;
            16'd12769: data <= 8'h07;
            16'd12770: data <= 8'hE0;
            16'd12771: data <= 8'h07;
            16'd12772: data <= 8'hE0;
            16'd12773: data <= 8'h07;
            16'd12774: data <= 8'hE0;
            16'd12775: data <= 8'h07;
            16'd12776: data <= 8'hE0;
            16'd12777: data <= 8'h07;
            16'd12778: data <= 8'hE0;
            16'd12779: data <= 8'h07;
            16'd12780: data <= 8'hE0;
            16'd12781: data <= 8'h07;
            16'd12782: data <= 8'hE0;
            16'd12783: data <= 8'h07;
            16'd12784: data <= 8'hE0;
            16'd12785: data <= 8'h07;
            16'd12786: data <= 8'hE0;
            16'd12787: data <= 8'h07;
            16'd12788: data <= 8'hE0;
            16'd12789: data <= 8'h07;
            16'd12790: data <= 8'hE0;
            16'd12791: data <= 8'h07;
            16'd12792: data <= 8'hE0;
            16'd12793: data <= 8'h07;
            16'd12794: data <= 8'hE0;
            16'd12795: data <= 8'h07;
            16'd12796: data <= 8'hE0;
            16'd12797: data <= 8'h07;
            16'd12798: data <= 8'hE0;
            16'd12799: data <= 8'h07;
            16'd12800: data <= 8'hFF;
            16'd12801: data <= 8'hFF;
            16'd12802: data <= 8'hE0;
            16'd12803: data <= 8'h07;
            16'd12804: data <= 8'hE0;
            16'd12805: data <= 8'h07;
            16'd12806: data <= 8'hE0;
            16'd12807: data <= 8'h07;
            16'd12808: data <= 8'hE0;
            16'd12809: data <= 8'h07;
            16'd12810: data <= 8'hE0;
            16'd12811: data <= 8'h07;
            16'd12812: data <= 8'hE0;
            16'd12813: data <= 8'h07;
            16'd12814: data <= 8'hE0;
            16'd12815: data <= 8'h07;
            16'd12816: data <= 8'hE0;
            16'd12817: data <= 8'h07;
            16'd12818: data <= 8'hE0;
            16'd12819: data <= 8'h07;
            16'd12820: data <= 8'hE0;
            16'd12821: data <= 8'h07;
            16'd12822: data <= 8'hE0;
            16'd12823: data <= 8'h07;
            16'd12824: data <= 8'hE0;
            16'd12825: data <= 8'h07;
            16'd12826: data <= 8'hE0;
            16'd12827: data <= 8'h07;
            16'd12828: data <= 8'hE0;
            16'd12829: data <= 8'h07;
            16'd12830: data <= 8'hE0;
            16'd12831: data <= 8'h07;
            16'd12832: data <= 8'hE0;
            16'd12833: data <= 8'h07;
            16'd12834: data <= 8'hE0;
            16'd12835: data <= 8'h07;
            16'd12836: data <= 8'hE0;
            16'd12837: data <= 8'h07;
            16'd12838: data <= 8'hE0;
            16'd12839: data <= 8'h07;
            16'd12840: data <= 8'hFF;
            16'd12841: data <= 8'hFF;
            16'd12842: data <= 8'hE0;
            16'd12843: data <= 8'h07;
            16'd12844: data <= 8'hE0;
            16'd12845: data <= 8'h07;
            16'd12846: data <= 8'hE0;
            16'd12847: data <= 8'h07;
            16'd12848: data <= 8'hE0;
            16'd12849: data <= 8'h07;
            16'd12850: data <= 8'hE0;
            16'd12851: data <= 8'h07;
            16'd12852: data <= 8'hE0;
            16'd12853: data <= 8'h07;
            16'd12854: data <= 8'hE0;
            16'd12855: data <= 8'h07;
            16'd12856: data <= 8'hE0;
            16'd12857: data <= 8'h07;
            16'd12858: data <= 8'hE0;
            16'd12859: data <= 8'h07;
            16'd12860: data <= 8'hE0;
            16'd12861: data <= 8'h07;
            16'd12862: data <= 8'hE0;
            16'd12863: data <= 8'h07;
            16'd12864: data <= 8'hE0;
            16'd12865: data <= 8'h07;
            16'd12866: data <= 8'hE0;
            16'd12867: data <= 8'h07;
            16'd12868: data <= 8'hE0;
            16'd12869: data <= 8'h07;
            16'd12870: data <= 8'hE0;
            16'd12871: data <= 8'h07;
            16'd12872: data <= 8'hE0;
            16'd12873: data <= 8'h07;
            16'd12874: data <= 8'hE0;
            16'd12875: data <= 8'h07;
            16'd12876: data <= 8'hE0;
            16'd12877: data <= 8'h07;
            16'd12878: data <= 8'hE0;
            16'd12879: data <= 8'h07;
            16'd12880: data <= 8'hFF;
            16'd12881: data <= 8'hFF;
            16'd12882: data <= 8'hE0;
            16'd12883: data <= 8'h07;
            16'd12884: data <= 8'hE0;
            16'd12885: data <= 8'h07;
            16'd12886: data <= 8'hE0;
            16'd12887: data <= 8'h07;
            16'd12888: data <= 8'hE0;
            16'd12889: data <= 8'h07;
            16'd12890: data <= 8'hE0;
            16'd12891: data <= 8'h07;
            16'd12892: data <= 8'hE0;
            16'd12893: data <= 8'h07;
            16'd12894: data <= 8'hE0;
            16'd12895: data <= 8'h07;
            16'd12896: data <= 8'hE0;
            16'd12897: data <= 8'h07;
            16'd12898: data <= 8'hE0;
            16'd12899: data <= 8'h07;
            16'd12900: data <= 8'hE0;
            16'd12901: data <= 8'h07;
            16'd12902: data <= 8'hE0;
            16'd12903: data <= 8'h07;
            16'd12904: data <= 8'hE0;
            16'd12905: data <= 8'h07;
            16'd12906: data <= 8'hE0;
            16'd12907: data <= 8'h07;
            16'd12908: data <= 8'hE0;
            16'd12909: data <= 8'h07;
            16'd12910: data <= 8'hE0;
            16'd12911: data <= 8'h07;
            16'd12912: data <= 8'hE0;
            16'd12913: data <= 8'h07;
            16'd12914: data <= 8'hE0;
            16'd12915: data <= 8'h07;
            16'd12916: data <= 8'hE0;
            16'd12917: data <= 8'h07;
            16'd12918: data <= 8'hE0;
            16'd12919: data <= 8'h07;
            16'd12920: data <= 8'hFF;
            16'd12921: data <= 8'hFF;
            16'd12922: data <= 8'hE0;
            16'd12923: data <= 8'h07;
            16'd12924: data <= 8'hE0;
            16'd12925: data <= 8'h07;
            16'd12926: data <= 8'hE0;
            16'd12927: data <= 8'h07;
            16'd12928: data <= 8'hE0;
            16'd12929: data <= 8'h07;
            16'd12930: data <= 8'hE0;
            16'd12931: data <= 8'h07;
            16'd12932: data <= 8'hE0;
            16'd12933: data <= 8'h07;
            16'd12934: data <= 8'hE0;
            16'd12935: data <= 8'h07;
            16'd12936: data <= 8'hE0;
            16'd12937: data <= 8'h07;
            16'd12938: data <= 8'hE0;
            16'd12939: data <= 8'h07;
            16'd12940: data <= 8'hE0;
            16'd12941: data <= 8'h07;
            16'd12942: data <= 8'hE0;
            16'd12943: data <= 8'h07;
            16'd12944: data <= 8'hE0;
            16'd12945: data <= 8'h07;
            16'd12946: data <= 8'hE0;
            16'd12947: data <= 8'h07;
            16'd12948: data <= 8'hE0;
            16'd12949: data <= 8'h07;
            16'd12950: data <= 8'hE0;
            16'd12951: data <= 8'h07;
            16'd12952: data <= 8'hE0;
            16'd12953: data <= 8'h07;
            16'd12954: data <= 8'hE0;
            16'd12955: data <= 8'h07;
            16'd12956: data <= 8'hE0;
            16'd12957: data <= 8'h07;
            16'd12958: data <= 8'hE0;
            16'd12959: data <= 8'h07;
            16'd12960: data <= 8'hFF;
            16'd12961: data <= 8'hFF;
            16'd12962: data <= 8'hE0;
            16'd12963: data <= 8'h07;
            16'd12964: data <= 8'hE0;
            16'd12965: data <= 8'h07;
            16'd12966: data <= 8'hE0;
            16'd12967: data <= 8'h07;
            16'd12968: data <= 8'hE0;
            16'd12969: data <= 8'h07;
            16'd12970: data <= 8'hE0;
            16'd12971: data <= 8'h07;
            16'd12972: data <= 8'hE0;
            16'd12973: data <= 8'h07;
            16'd12974: data <= 8'hE0;
            16'd12975: data <= 8'h07;
            16'd12976: data <= 8'hE0;
            16'd12977: data <= 8'h07;
            16'd12978: data <= 8'hE0;
            16'd12979: data <= 8'h07;
            16'd12980: data <= 8'hE0;
            16'd12981: data <= 8'h07;
            16'd12982: data <= 8'hE0;
            16'd12983: data <= 8'h07;
            16'd12984: data <= 8'hE0;
            16'd12985: data <= 8'h07;
            16'd12986: data <= 8'hE0;
            16'd12987: data <= 8'h07;
            16'd12988: data <= 8'hE0;
            16'd12989: data <= 8'h07;
            16'd12990: data <= 8'hE0;
            16'd12991: data <= 8'h07;
            16'd12992: data <= 8'hE0;
            16'd12993: data <= 8'h07;
            16'd12994: data <= 8'hE0;
            16'd12995: data <= 8'h07;
            16'd12996: data <= 8'hE0;
            16'd12997: data <= 8'h07;
            16'd12998: data <= 8'hE0;
            16'd12999: data <= 8'h07;
            16'd13000: data <= 8'hFF;
            16'd13001: data <= 8'hFF;
            16'd13002: data <= 8'hE0;
            16'd13003: data <= 8'h07;
            16'd13004: data <= 8'hE0;
            16'd13005: data <= 8'h07;
            16'd13006: data <= 8'hE0;
            16'd13007: data <= 8'h07;
            16'd13008: data <= 8'hE0;
            16'd13009: data <= 8'h07;
            16'd13010: data <= 8'hE0;
            16'd13011: data <= 8'h07;
            16'd13012: data <= 8'hE0;
            16'd13013: data <= 8'h07;
            16'd13014: data <= 8'hE0;
            16'd13015: data <= 8'h07;
            16'd13016: data <= 8'hE0;
            16'd13017: data <= 8'h07;
            16'd13018: data <= 8'hE0;
            16'd13019: data <= 8'h07;
            16'd13020: data <= 8'hE0;
            16'd13021: data <= 8'h07;
            16'd13022: data <= 8'hE0;
            16'd13023: data <= 8'h07;
            16'd13024: data <= 8'hE0;
            16'd13025: data <= 8'h07;
            16'd13026: data <= 8'hE0;
            16'd13027: data <= 8'h07;
            16'd13028: data <= 8'hE0;
            16'd13029: data <= 8'h07;
            16'd13030: data <= 8'hE0;
            16'd13031: data <= 8'h07;
            16'd13032: data <= 8'hE0;
            16'd13033: data <= 8'h07;
            16'd13034: data <= 8'hE0;
            16'd13035: data <= 8'h07;
            16'd13036: data <= 8'hE0;
            16'd13037: data <= 8'h07;
            16'd13038: data <= 8'hE0;
            16'd13039: data <= 8'h07;
            16'd13040: data <= 8'hFF;
            16'd13041: data <= 8'hFF;
            16'd13042: data <= 8'hE0;
            16'd13043: data <= 8'h07;
            16'd13044: data <= 8'hE0;
            16'd13045: data <= 8'h07;
            16'd13046: data <= 8'hE0;
            16'd13047: data <= 8'h07;
            16'd13048: data <= 8'hE0;
            16'd13049: data <= 8'h07;
            16'd13050: data <= 8'hE0;
            16'd13051: data <= 8'h07;
            16'd13052: data <= 8'hE0;
            16'd13053: data <= 8'h07;
            16'd13054: data <= 8'hE0;
            16'd13055: data <= 8'h07;
            16'd13056: data <= 8'hE0;
            16'd13057: data <= 8'h07;
            16'd13058: data <= 8'hE0;
            16'd13059: data <= 8'h07;
            16'd13060: data <= 8'hE0;
            16'd13061: data <= 8'h07;
            16'd13062: data <= 8'hE0;
            16'd13063: data <= 8'h07;
            16'd13064: data <= 8'hE0;
            16'd13065: data <= 8'h07;
            16'd13066: data <= 8'hE0;
            16'd13067: data <= 8'h07;
            16'd13068: data <= 8'hE0;
            16'd13069: data <= 8'h07;
            16'd13070: data <= 8'hE0;
            16'd13071: data <= 8'h07;
            16'd13072: data <= 8'hE0;
            16'd13073: data <= 8'h07;
            16'd13074: data <= 8'hE0;
            16'd13075: data <= 8'h07;
            16'd13076: data <= 8'hE0;
            16'd13077: data <= 8'h07;
            16'd13078: data <= 8'hE0;
            16'd13079: data <= 8'h07;
            16'd13080: data <= 8'hFF;
            16'd13081: data <= 8'hFF;
            16'd13082: data <= 8'hE0;
            16'd13083: data <= 8'h07;
            16'd13084: data <= 8'hE0;
            16'd13085: data <= 8'h07;
            16'd13086: data <= 8'hE0;
            16'd13087: data <= 8'h07;
            16'd13088: data <= 8'hE0;
            16'd13089: data <= 8'h07;
            16'd13090: data <= 8'hE0;
            16'd13091: data <= 8'h07;
            16'd13092: data <= 8'hE0;
            16'd13093: data <= 8'h07;
            16'd13094: data <= 8'hE0;
            16'd13095: data <= 8'h07;
            16'd13096: data <= 8'hE0;
            16'd13097: data <= 8'h07;
            16'd13098: data <= 8'hE0;
            16'd13099: data <= 8'h07;
            16'd13100: data <= 8'hE0;
            16'd13101: data <= 8'h07;
            16'd13102: data <= 8'hE0;
            16'd13103: data <= 8'h07;
            16'd13104: data <= 8'hE0;
            16'd13105: data <= 8'h07;
            16'd13106: data <= 8'hE0;
            16'd13107: data <= 8'h07;
            16'd13108: data <= 8'hE0;
            16'd13109: data <= 8'h07;
            16'd13110: data <= 8'hE0;
            16'd13111: data <= 8'h07;
            16'd13112: data <= 8'hE0;
            16'd13113: data <= 8'h07;
            16'd13114: data <= 8'hE0;
            16'd13115: data <= 8'h07;
            16'd13116: data <= 8'hE0;
            16'd13117: data <= 8'h07;
            16'd13118: data <= 8'hE0;
            16'd13119: data <= 8'h07;
            16'd13120: data <= 8'hFF;
            16'd13121: data <= 8'hFF;
            16'd13122: data <= 8'hE0;
            16'd13123: data <= 8'h07;
            16'd13124: data <= 8'hE0;
            16'd13125: data <= 8'h07;
            16'd13126: data <= 8'hE0;
            16'd13127: data <= 8'h07;
            16'd13128: data <= 8'hE0;
            16'd13129: data <= 8'h07;
            16'd13130: data <= 8'hE0;
            16'd13131: data <= 8'h07;
            16'd13132: data <= 8'hE0;
            16'd13133: data <= 8'h07;
            16'd13134: data <= 8'hE0;
            16'd13135: data <= 8'h07;
            16'd13136: data <= 8'hE0;
            16'd13137: data <= 8'h07;
            16'd13138: data <= 8'hE0;
            16'd13139: data <= 8'h07;
            16'd13140: data <= 8'hE0;
            16'd13141: data <= 8'h07;
            16'd13142: data <= 8'hE0;
            16'd13143: data <= 8'h07;
            16'd13144: data <= 8'hE0;
            16'd13145: data <= 8'h07;
            16'd13146: data <= 8'hE0;
            16'd13147: data <= 8'h07;
            16'd13148: data <= 8'hE0;
            16'd13149: data <= 8'h07;
            16'd13150: data <= 8'hE0;
            16'd13151: data <= 8'h07;
            16'd13152: data <= 8'hE0;
            16'd13153: data <= 8'h07;
            16'd13154: data <= 8'hE0;
            16'd13155: data <= 8'h07;
            16'd13156: data <= 8'hE0;
            16'd13157: data <= 8'h07;
            16'd13158: data <= 8'hE0;
            16'd13159: data <= 8'h07;
            16'd13160: data <= 8'hFF;
            16'd13161: data <= 8'hFF;
            16'd13162: data <= 8'hE0;
            16'd13163: data <= 8'h07;
            16'd13164: data <= 8'hE0;
            16'd13165: data <= 8'h07;
            16'd13166: data <= 8'hE0;
            16'd13167: data <= 8'h07;
            16'd13168: data <= 8'hE0;
            16'd13169: data <= 8'h07;
            16'd13170: data <= 8'hE0;
            16'd13171: data <= 8'h07;
            16'd13172: data <= 8'hE0;
            16'd13173: data <= 8'h07;
            16'd13174: data <= 8'hE0;
            16'd13175: data <= 8'h07;
            16'd13176: data <= 8'hE0;
            16'd13177: data <= 8'h07;
            16'd13178: data <= 8'hE0;
            16'd13179: data <= 8'h07;
            16'd13180: data <= 8'hE0;
            16'd13181: data <= 8'h07;
            16'd13182: data <= 8'hE0;
            16'd13183: data <= 8'h07;
            16'd13184: data <= 8'hE0;
            16'd13185: data <= 8'h07;
            16'd13186: data <= 8'hE0;
            16'd13187: data <= 8'h07;
            16'd13188: data <= 8'hE0;
            16'd13189: data <= 8'h07;
            16'd13190: data <= 8'hE0;
            16'd13191: data <= 8'h07;
            16'd13192: data <= 8'hE0;
            16'd13193: data <= 8'h07;
            16'd13194: data <= 8'hE0;
            16'd13195: data <= 8'h07;
            16'd13196: data <= 8'hE0;
            16'd13197: data <= 8'h07;
            16'd13198: data <= 8'hE0;
            16'd13199: data <= 8'h07;
            16'd13200: data <= 8'hFF;
            16'd13201: data <= 8'hFF;
            16'd13202: data <= 8'hE0;
            16'd13203: data <= 8'h07;
            16'd13204: data <= 8'hE0;
            16'd13205: data <= 8'h07;
            16'd13206: data <= 8'hE0;
            16'd13207: data <= 8'h07;
            16'd13208: data <= 8'hE0;
            16'd13209: data <= 8'h07;
            16'd13210: data <= 8'hE0;
            16'd13211: data <= 8'h07;
            16'd13212: data <= 8'hE0;
            16'd13213: data <= 8'h07;
            16'd13214: data <= 8'hE0;
            16'd13215: data <= 8'h07;
            16'd13216: data <= 8'hE0;
            16'd13217: data <= 8'h07;
            16'd13218: data <= 8'hE0;
            16'd13219: data <= 8'h07;
            16'd13220: data <= 8'hE0;
            16'd13221: data <= 8'h07;
            16'd13222: data <= 8'hE0;
            16'd13223: data <= 8'h07;
            16'd13224: data <= 8'hE0;
            16'd13225: data <= 8'h07;
            16'd13226: data <= 8'hE0;
            16'd13227: data <= 8'h07;
            16'd13228: data <= 8'hE0;
            16'd13229: data <= 8'h07;
            16'd13230: data <= 8'hE0;
            16'd13231: data <= 8'h07;
            16'd13232: data <= 8'hE0;
            16'd13233: data <= 8'h07;
            16'd13234: data <= 8'hE0;
            16'd13235: data <= 8'h07;
            16'd13236: data <= 8'hE0;
            16'd13237: data <= 8'h07;
            16'd13238: data <= 8'hE0;
            16'd13239: data <= 8'h07;
            16'd13240: data <= 8'hFF;
            16'd13241: data <= 8'hFF;
            16'd13242: data <= 8'hE0;
            16'd13243: data <= 8'h07;
            16'd13244: data <= 8'hE0;
            16'd13245: data <= 8'h07;
            16'd13246: data <= 8'hE0;
            16'd13247: data <= 8'h07;
            16'd13248: data <= 8'hE0;
            16'd13249: data <= 8'h07;
            16'd13250: data <= 8'hE0;
            16'd13251: data <= 8'h07;
            16'd13252: data <= 8'hE0;
            16'd13253: data <= 8'h07;
            16'd13254: data <= 8'hE0;
            16'd13255: data <= 8'h07;
            16'd13256: data <= 8'hE0;
            16'd13257: data <= 8'h07;
            16'd13258: data <= 8'hE0;
            16'd13259: data <= 8'h07;
            16'd13260: data <= 8'hE0;
            16'd13261: data <= 8'h07;
            16'd13262: data <= 8'hE0;
            16'd13263: data <= 8'h07;
            16'd13264: data <= 8'hE0;
            16'd13265: data <= 8'h07;
            16'd13266: data <= 8'hE0;
            16'd13267: data <= 8'h07;
            16'd13268: data <= 8'hE0;
            16'd13269: data <= 8'h07;
            16'd13270: data <= 8'hE0;
            16'd13271: data <= 8'h07;
            16'd13272: data <= 8'hE0;
            16'd13273: data <= 8'h07;
            16'd13274: data <= 8'hE0;
            16'd13275: data <= 8'h07;
            16'd13276: data <= 8'hE0;
            16'd13277: data <= 8'h07;
            16'd13278: data <= 8'hE0;
            16'd13279: data <= 8'h07;
            16'd13280: data <= 8'hFF;
            16'd13281: data <= 8'hFF;
            16'd13282: data <= 8'hE0;
            16'd13283: data <= 8'h07;
            16'd13284: data <= 8'hE0;
            16'd13285: data <= 8'h07;
            16'd13286: data <= 8'hE0;
            16'd13287: data <= 8'h07;
            16'd13288: data <= 8'hE0;
            16'd13289: data <= 8'h07;
            16'd13290: data <= 8'hE0;
            16'd13291: data <= 8'h07;
            16'd13292: data <= 8'hE0;
            16'd13293: data <= 8'h07;
            16'd13294: data <= 8'hE0;
            16'd13295: data <= 8'h07;
            16'd13296: data <= 8'hE0;
            16'd13297: data <= 8'h07;
            16'd13298: data <= 8'hE0;
            16'd13299: data <= 8'h07;
            16'd13300: data <= 8'hE0;
            16'd13301: data <= 8'h07;
            16'd13302: data <= 8'hE0;
            16'd13303: data <= 8'h07;
            16'd13304: data <= 8'hE0;
            16'd13305: data <= 8'h07;
            16'd13306: data <= 8'hE0;
            16'd13307: data <= 8'h07;
            16'd13308: data <= 8'hE0;
            16'd13309: data <= 8'h07;
            16'd13310: data <= 8'hE0;
            16'd13311: data <= 8'h07;
            16'd13312: data <= 8'hE0;
            16'd13313: data <= 8'h07;
            16'd13314: data <= 8'hE0;
            16'd13315: data <= 8'h07;
            16'd13316: data <= 8'hE0;
            16'd13317: data <= 8'h07;
            16'd13318: data <= 8'hE0;
            16'd13319: data <= 8'h07;
            16'd13320: data <= 8'hFF;
            16'd13321: data <= 8'hFF;
            16'd13322: data <= 8'hE0;
            16'd13323: data <= 8'h07;
            16'd13324: data <= 8'hE0;
            16'd13325: data <= 8'h07;
            16'd13326: data <= 8'hE0;
            16'd13327: data <= 8'h07;
            16'd13328: data <= 8'hE0;
            16'd13329: data <= 8'h07;
            16'd13330: data <= 8'hE0;
            16'd13331: data <= 8'h07;
            16'd13332: data <= 8'hE0;
            16'd13333: data <= 8'h07;
            16'd13334: data <= 8'hE0;
            16'd13335: data <= 8'h07;
            16'd13336: data <= 8'hE0;
            16'd13337: data <= 8'h07;
            16'd13338: data <= 8'hE0;
            16'd13339: data <= 8'h07;
            16'd13340: data <= 8'hE0;
            16'd13341: data <= 8'h07;
            16'd13342: data <= 8'hE0;
            16'd13343: data <= 8'h07;
            16'd13344: data <= 8'hE0;
            16'd13345: data <= 8'h07;
            16'd13346: data <= 8'hE0;
            16'd13347: data <= 8'h07;
            16'd13348: data <= 8'hE0;
            16'd13349: data <= 8'h07;
            16'd13350: data <= 8'hE0;
            16'd13351: data <= 8'h07;
            16'd13352: data <= 8'hE0;
            16'd13353: data <= 8'h07;
            16'd13354: data <= 8'hE0;
            16'd13355: data <= 8'h07;
            16'd13356: data <= 8'hE0;
            16'd13357: data <= 8'h07;
            16'd13358: data <= 8'hE0;
            16'd13359: data <= 8'h07;
            16'd13360: data <= 8'hFF;
            16'd13361: data <= 8'hFF;
            16'd13362: data <= 8'hE0;
            16'd13363: data <= 8'h07;
            16'd13364: data <= 8'hE0;
            16'd13365: data <= 8'h07;
            16'd13366: data <= 8'hE0;
            16'd13367: data <= 8'h07;
            16'd13368: data <= 8'hE0;
            16'd13369: data <= 8'h07;
            16'd13370: data <= 8'hE0;
            16'd13371: data <= 8'h07;
            16'd13372: data <= 8'hE0;
            16'd13373: data <= 8'h07;
            16'd13374: data <= 8'hE0;
            16'd13375: data <= 8'h07;
            16'd13376: data <= 8'hE0;
            16'd13377: data <= 8'h07;
            16'd13378: data <= 8'hE0;
            16'd13379: data <= 8'h07;
            16'd13380: data <= 8'hE0;
            16'd13381: data <= 8'h07;
            16'd13382: data <= 8'hE0;
            16'd13383: data <= 8'h07;
            16'd13384: data <= 8'hE0;
            16'd13385: data <= 8'h07;
            16'd13386: data <= 8'hE0;
            16'd13387: data <= 8'h07;
            16'd13388: data <= 8'hE0;
            16'd13389: data <= 8'h07;
            16'd13390: data <= 8'hE0;
            16'd13391: data <= 8'h07;
            16'd13392: data <= 8'hE0;
            16'd13393: data <= 8'h07;
            16'd13394: data <= 8'hE0;
            16'd13395: data <= 8'h07;
            16'd13396: data <= 8'hE0;
            16'd13397: data <= 8'h07;
            16'd13398: data <= 8'hE0;
            16'd13399: data <= 8'h07;
            16'd13400: data <= 8'hFF;
            16'd13401: data <= 8'hFF;
            16'd13402: data <= 8'hE0;
            16'd13403: data <= 8'h07;
            16'd13404: data <= 8'hE0;
            16'd13405: data <= 8'h07;
            16'd13406: data <= 8'hE0;
            16'd13407: data <= 8'h07;
            16'd13408: data <= 8'hE0;
            16'd13409: data <= 8'h07;
            16'd13410: data <= 8'hE0;
            16'd13411: data <= 8'h07;
            16'd13412: data <= 8'hE0;
            16'd13413: data <= 8'h07;
            16'd13414: data <= 8'hE0;
            16'd13415: data <= 8'h07;
            16'd13416: data <= 8'hE0;
            16'd13417: data <= 8'h07;
            16'd13418: data <= 8'hE0;
            16'd13419: data <= 8'h07;
            16'd13420: data <= 8'hE0;
            16'd13421: data <= 8'h07;
            16'd13422: data <= 8'hE0;
            16'd13423: data <= 8'h07;
            16'd13424: data <= 8'hE0;
            16'd13425: data <= 8'h07;
            16'd13426: data <= 8'hE0;
            16'd13427: data <= 8'h07;
            16'd13428: data <= 8'hE0;
            16'd13429: data <= 8'h07;
            16'd13430: data <= 8'hE0;
            16'd13431: data <= 8'h07;
            16'd13432: data <= 8'hE0;
            16'd13433: data <= 8'h07;
            16'd13434: data <= 8'hE0;
            16'd13435: data <= 8'h07;
            16'd13436: data <= 8'hE0;
            16'd13437: data <= 8'h07;
            16'd13438: data <= 8'hE0;
            16'd13439: data <= 8'h07;
            16'd13440: data <= 8'hFF;
            16'd13441: data <= 8'hFF;
            16'd13442: data <= 8'hE0;
            16'd13443: data <= 8'h07;
            16'd13444: data <= 8'hE0;
            16'd13445: data <= 8'h07;
            16'd13446: data <= 8'hE0;
            16'd13447: data <= 8'h07;
            16'd13448: data <= 8'hE0;
            16'd13449: data <= 8'h07;
            16'd13450: data <= 8'hE0;
            16'd13451: data <= 8'h07;
            16'd13452: data <= 8'hE0;
            16'd13453: data <= 8'h07;
            16'd13454: data <= 8'hE0;
            16'd13455: data <= 8'h07;
            16'd13456: data <= 8'hE0;
            16'd13457: data <= 8'h07;
            16'd13458: data <= 8'hE0;
            16'd13459: data <= 8'h07;
            16'd13460: data <= 8'hE0;
            16'd13461: data <= 8'h07;
            16'd13462: data <= 8'hE0;
            16'd13463: data <= 8'h07;
            16'd13464: data <= 8'hE0;
            16'd13465: data <= 8'h07;
            16'd13466: data <= 8'hE0;
            16'd13467: data <= 8'h07;
            16'd13468: data <= 8'hE0;
            16'd13469: data <= 8'h07;
            16'd13470: data <= 8'hE0;
            16'd13471: data <= 8'h07;
            16'd13472: data <= 8'hE0;
            16'd13473: data <= 8'h07;
            16'd13474: data <= 8'hE0;
            16'd13475: data <= 8'h07;
            16'd13476: data <= 8'hE0;
            16'd13477: data <= 8'h07;
            16'd13478: data <= 8'hE0;
            16'd13479: data <= 8'h07;
            16'd13480: data <= 8'hFF;
            16'd13481: data <= 8'hFF;
            16'd13482: data <= 8'hE0;
            16'd13483: data <= 8'h07;
            16'd13484: data <= 8'hE0;
            16'd13485: data <= 8'h07;
            16'd13486: data <= 8'hE0;
            16'd13487: data <= 8'h07;
            16'd13488: data <= 8'hE0;
            16'd13489: data <= 8'h07;
            16'd13490: data <= 8'hE0;
            16'd13491: data <= 8'h07;
            16'd13492: data <= 8'hE0;
            16'd13493: data <= 8'h07;
            16'd13494: data <= 8'hE0;
            16'd13495: data <= 8'h07;
            16'd13496: data <= 8'hE0;
            16'd13497: data <= 8'h07;
            16'd13498: data <= 8'hE0;
            16'd13499: data <= 8'h07;
            16'd13500: data <= 8'hE0;
            16'd13501: data <= 8'h07;
            16'd13502: data <= 8'hE0;
            16'd13503: data <= 8'h07;
            16'd13504: data <= 8'hE0;
            16'd13505: data <= 8'h07;
            16'd13506: data <= 8'hE0;
            16'd13507: data <= 8'h07;
            16'd13508: data <= 8'hE0;
            16'd13509: data <= 8'h07;
            16'd13510: data <= 8'hE0;
            16'd13511: data <= 8'h07;
            16'd13512: data <= 8'hE0;
            16'd13513: data <= 8'h07;
            16'd13514: data <= 8'hE0;
            16'd13515: data <= 8'h07;
            16'd13516: data <= 8'hE0;
            16'd13517: data <= 8'h07;
            16'd13518: data <= 8'hE0;
            16'd13519: data <= 8'h07;
            16'd13520: data <= 8'hFF;
            16'd13521: data <= 8'hFF;
            16'd13522: data <= 8'hE0;
            16'd13523: data <= 8'h07;
            16'd13524: data <= 8'hE0;
            16'd13525: data <= 8'h07;
            16'd13526: data <= 8'hE0;
            16'd13527: data <= 8'h07;
            16'd13528: data <= 8'hE0;
            16'd13529: data <= 8'h07;
            16'd13530: data <= 8'hE0;
            16'd13531: data <= 8'h07;
            16'd13532: data <= 8'hE0;
            16'd13533: data <= 8'h07;
            16'd13534: data <= 8'hE0;
            16'd13535: data <= 8'h07;
            16'd13536: data <= 8'hE0;
            16'd13537: data <= 8'h07;
            16'd13538: data <= 8'hE0;
            16'd13539: data <= 8'h07;
            16'd13540: data <= 8'hE0;
            16'd13541: data <= 8'h07;
            16'd13542: data <= 8'hE0;
            16'd13543: data <= 8'h07;
            16'd13544: data <= 8'hE0;
            16'd13545: data <= 8'h07;
            16'd13546: data <= 8'hE0;
            16'd13547: data <= 8'h07;
            16'd13548: data <= 8'hE0;
            16'd13549: data <= 8'h07;
            16'd13550: data <= 8'hE0;
            16'd13551: data <= 8'h07;
            16'd13552: data <= 8'hE0;
            16'd13553: data <= 8'h07;
            16'd13554: data <= 8'hE0;
            16'd13555: data <= 8'h07;
            16'd13556: data <= 8'hE0;
            16'd13557: data <= 8'h07;
            16'd13558: data <= 8'hE0;
            16'd13559: data <= 8'h07;
            16'd13560: data <= 8'hFF;
            16'd13561: data <= 8'hFF;
            16'd13562: data <= 8'hE0;
            16'd13563: data <= 8'h07;
            16'd13564: data <= 8'hE0;
            16'd13565: data <= 8'h07;
            16'd13566: data <= 8'hE0;
            16'd13567: data <= 8'h07;
            16'd13568: data <= 8'hE0;
            16'd13569: data <= 8'h07;
            16'd13570: data <= 8'hE0;
            16'd13571: data <= 8'h07;
            16'd13572: data <= 8'hE0;
            16'd13573: data <= 8'h07;
            16'd13574: data <= 8'hE0;
            16'd13575: data <= 8'h07;
            16'd13576: data <= 8'hE0;
            16'd13577: data <= 8'h07;
            16'd13578: data <= 8'hE0;
            16'd13579: data <= 8'h07;
            16'd13580: data <= 8'hE0;
            16'd13581: data <= 8'h07;
            16'd13582: data <= 8'hE0;
            16'd13583: data <= 8'h07;
            16'd13584: data <= 8'hE0;
            16'd13585: data <= 8'h07;
            16'd13586: data <= 8'hE0;
            16'd13587: data <= 8'h07;
            16'd13588: data <= 8'hE0;
            16'd13589: data <= 8'h07;
            16'd13590: data <= 8'hE0;
            16'd13591: data <= 8'h07;
            16'd13592: data <= 8'hE0;
            16'd13593: data <= 8'h07;
            16'd13594: data <= 8'hE0;
            16'd13595: data <= 8'h07;
            16'd13596: data <= 8'hE0;
            16'd13597: data <= 8'h07;
            16'd13598: data <= 8'hE0;
            16'd13599: data <= 8'h07;
            16'd13600: data <= 8'hFF;
            16'd13601: data <= 8'hFF;
            16'd13602: data <= 8'hE0;
            16'd13603: data <= 8'h07;
            16'd13604: data <= 8'hE0;
            16'd13605: data <= 8'h07;
            16'd13606: data <= 8'hE0;
            16'd13607: data <= 8'h07;
            16'd13608: data <= 8'hE0;
            16'd13609: data <= 8'h07;
            16'd13610: data <= 8'hE0;
            16'd13611: data <= 8'h07;
            16'd13612: data <= 8'hE0;
            16'd13613: data <= 8'h07;
            16'd13614: data <= 8'hE0;
            16'd13615: data <= 8'h07;
            16'd13616: data <= 8'hE0;
            16'd13617: data <= 8'h07;
            16'd13618: data <= 8'hE0;
            16'd13619: data <= 8'h07;
            16'd13620: data <= 8'hE0;
            16'd13621: data <= 8'h07;
            16'd13622: data <= 8'hE0;
            16'd13623: data <= 8'h07;
            16'd13624: data <= 8'hE0;
            16'd13625: data <= 8'h07;
            16'd13626: data <= 8'hE0;
            16'd13627: data <= 8'h07;
            16'd13628: data <= 8'hE0;
            16'd13629: data <= 8'h07;
            16'd13630: data <= 8'hE0;
            16'd13631: data <= 8'h07;
            16'd13632: data <= 8'hE0;
            16'd13633: data <= 8'h07;
            16'd13634: data <= 8'hE0;
            16'd13635: data <= 8'h07;
            16'd13636: data <= 8'hE0;
            16'd13637: data <= 8'h07;
            16'd13638: data <= 8'hE0;
            16'd13639: data <= 8'h07;
            16'd13640: data <= 8'hFF;
            16'd13641: data <= 8'hFF;
            16'd13642: data <= 8'hE0;
            16'd13643: data <= 8'h07;
            16'd13644: data <= 8'hE0;
            16'd13645: data <= 8'h07;
            16'd13646: data <= 8'hE0;
            16'd13647: data <= 8'h07;
            16'd13648: data <= 8'hE0;
            16'd13649: data <= 8'h07;
            16'd13650: data <= 8'hE0;
            16'd13651: data <= 8'h07;
            16'd13652: data <= 8'hE0;
            16'd13653: data <= 8'h07;
            16'd13654: data <= 8'hE0;
            16'd13655: data <= 8'h07;
            16'd13656: data <= 8'hE0;
            16'd13657: data <= 8'h07;
            16'd13658: data <= 8'hE0;
            16'd13659: data <= 8'h07;
            16'd13660: data <= 8'hE0;
            16'd13661: data <= 8'h07;
            16'd13662: data <= 8'hE0;
            16'd13663: data <= 8'h07;
            16'd13664: data <= 8'hE0;
            16'd13665: data <= 8'h07;
            16'd13666: data <= 8'hE0;
            16'd13667: data <= 8'h07;
            16'd13668: data <= 8'hE0;
            16'd13669: data <= 8'h07;
            16'd13670: data <= 8'hE0;
            16'd13671: data <= 8'h07;
            16'd13672: data <= 8'hE0;
            16'd13673: data <= 8'h07;
            16'd13674: data <= 8'hE0;
            16'd13675: data <= 8'h07;
            16'd13676: data <= 8'hE0;
            16'd13677: data <= 8'h07;
            16'd13678: data <= 8'hE0;
            16'd13679: data <= 8'h07;
            16'd13680: data <= 8'hFF;
            16'd13681: data <= 8'hFF;
            16'd13682: data <= 8'hE0;
            16'd13683: data <= 8'h07;
            16'd13684: data <= 8'hE0;
            16'd13685: data <= 8'h07;
            16'd13686: data <= 8'hE0;
            16'd13687: data <= 8'h07;
            16'd13688: data <= 8'hE0;
            16'd13689: data <= 8'h07;
            16'd13690: data <= 8'hE0;
            16'd13691: data <= 8'h07;
            16'd13692: data <= 8'hE0;
            16'd13693: data <= 8'h07;
            16'd13694: data <= 8'hE0;
            16'd13695: data <= 8'h07;
            16'd13696: data <= 8'hE0;
            16'd13697: data <= 8'h07;
            16'd13698: data <= 8'hE0;
            16'd13699: data <= 8'h07;
            16'd13700: data <= 8'hE0;
            16'd13701: data <= 8'h07;
            16'd13702: data <= 8'hE0;
            16'd13703: data <= 8'h07;
            16'd13704: data <= 8'hE0;
            16'd13705: data <= 8'h07;
            16'd13706: data <= 8'hE0;
            16'd13707: data <= 8'h07;
            16'd13708: data <= 8'hE0;
            16'd13709: data <= 8'h07;
            16'd13710: data <= 8'hE0;
            16'd13711: data <= 8'h07;
            16'd13712: data <= 8'hE0;
            16'd13713: data <= 8'h07;
            16'd13714: data <= 8'hE0;
            16'd13715: data <= 8'h07;
            16'd13716: data <= 8'hE0;
            16'd13717: data <= 8'h07;
            16'd13718: data <= 8'hE0;
            16'd13719: data <= 8'h07;
            16'd13720: data <= 8'hFF;
            16'd13721: data <= 8'hFF;
            16'd13722: data <= 8'hE0;
            16'd13723: data <= 8'h07;
            16'd13724: data <= 8'hE0;
            16'd13725: data <= 8'h07;
            16'd13726: data <= 8'hE0;
            16'd13727: data <= 8'h07;
            16'd13728: data <= 8'hE0;
            16'd13729: data <= 8'h07;
            16'd13730: data <= 8'hE0;
            16'd13731: data <= 8'h07;
            16'd13732: data <= 8'hE0;
            16'd13733: data <= 8'h07;
            16'd13734: data <= 8'hE0;
            16'd13735: data <= 8'h07;
            16'd13736: data <= 8'hE0;
            16'd13737: data <= 8'h07;
            16'd13738: data <= 8'hE0;
            16'd13739: data <= 8'h07;
            16'd13740: data <= 8'hE0;
            16'd13741: data <= 8'h07;
            16'd13742: data <= 8'hE0;
            16'd13743: data <= 8'h07;
            16'd13744: data <= 8'hE0;
            16'd13745: data <= 8'h07;
            16'd13746: data <= 8'hE0;
            16'd13747: data <= 8'h07;
            16'd13748: data <= 8'hE0;
            16'd13749: data <= 8'h07;
            16'd13750: data <= 8'hE0;
            16'd13751: data <= 8'h07;
            16'd13752: data <= 8'hE0;
            16'd13753: data <= 8'h07;
            16'd13754: data <= 8'hE0;
            16'd13755: data <= 8'h07;
            16'd13756: data <= 8'hE0;
            16'd13757: data <= 8'h07;
            16'd13758: data <= 8'hE0;
            16'd13759: data <= 8'h07;
            16'd13760: data <= 8'hFF;
            16'd13761: data <= 8'hFF;
            16'd13762: data <= 8'hE0;
            16'd13763: data <= 8'h07;
            16'd13764: data <= 8'hE0;
            16'd13765: data <= 8'h07;
            16'd13766: data <= 8'hE0;
            16'd13767: data <= 8'h07;
            16'd13768: data <= 8'hE0;
            16'd13769: data <= 8'h07;
            16'd13770: data <= 8'hE0;
            16'd13771: data <= 8'h07;
            16'd13772: data <= 8'hE0;
            16'd13773: data <= 8'h07;
            16'd13774: data <= 8'hE0;
            16'd13775: data <= 8'h07;
            16'd13776: data <= 8'hE0;
            16'd13777: data <= 8'h07;
            16'd13778: data <= 8'hE0;
            16'd13779: data <= 8'h07;
            16'd13780: data <= 8'hE0;
            16'd13781: data <= 8'h07;
            16'd13782: data <= 8'hE0;
            16'd13783: data <= 8'h07;
            16'd13784: data <= 8'hE0;
            16'd13785: data <= 8'h07;
            16'd13786: data <= 8'hE0;
            16'd13787: data <= 8'h07;
            16'd13788: data <= 8'hE0;
            16'd13789: data <= 8'h07;
            16'd13790: data <= 8'hE0;
            16'd13791: data <= 8'h07;
            16'd13792: data <= 8'hE0;
            16'd13793: data <= 8'h07;
            16'd13794: data <= 8'hE0;
            16'd13795: data <= 8'h07;
            16'd13796: data <= 8'hE0;
            16'd13797: data <= 8'h07;
            16'd13798: data <= 8'hE0;
            16'd13799: data <= 8'h07;
            16'd13800: data <= 8'hFF;
            16'd13801: data <= 8'hFF;
            16'd13802: data <= 8'hE0;
            16'd13803: data <= 8'h07;
            16'd13804: data <= 8'hE0;
            16'd13805: data <= 8'h07;
            16'd13806: data <= 8'hE0;
            16'd13807: data <= 8'h07;
            16'd13808: data <= 8'hE0;
            16'd13809: data <= 8'h07;
            16'd13810: data <= 8'hE0;
            16'd13811: data <= 8'h07;
            16'd13812: data <= 8'hE0;
            16'd13813: data <= 8'h07;
            16'd13814: data <= 8'hE0;
            16'd13815: data <= 8'h07;
            16'd13816: data <= 8'hE0;
            16'd13817: data <= 8'h07;
            16'd13818: data <= 8'hE0;
            16'd13819: data <= 8'h07;
            16'd13820: data <= 8'hE0;
            16'd13821: data <= 8'h07;
            16'd13822: data <= 8'hE0;
            16'd13823: data <= 8'h07;
            16'd13824: data <= 8'hE0;
            16'd13825: data <= 8'h07;
            16'd13826: data <= 8'hE0;
            16'd13827: data <= 8'h07;
            16'd13828: data <= 8'hE0;
            16'd13829: data <= 8'h07;
            16'd13830: data <= 8'hE0;
            16'd13831: data <= 8'h07;
            16'd13832: data <= 8'hE0;
            16'd13833: data <= 8'h07;
            16'd13834: data <= 8'hE0;
            16'd13835: data <= 8'h07;
            16'd13836: data <= 8'hE0;
            16'd13837: data <= 8'h07;
            16'd13838: data <= 8'hE0;
            16'd13839: data <= 8'h07;
            16'd13840: data <= 8'hFF;
            16'd13841: data <= 8'hFF;
            16'd13842: data <= 8'hE0;
            16'd13843: data <= 8'h07;
            16'd13844: data <= 8'hE0;
            16'd13845: data <= 8'h07;
            16'd13846: data <= 8'hE0;
            16'd13847: data <= 8'h07;
            16'd13848: data <= 8'hE0;
            16'd13849: data <= 8'h07;
            16'd13850: data <= 8'hE0;
            16'd13851: data <= 8'h07;
            16'd13852: data <= 8'hE0;
            16'd13853: data <= 8'h07;
            16'd13854: data <= 8'hE0;
            16'd13855: data <= 8'h07;
            16'd13856: data <= 8'hE0;
            16'd13857: data <= 8'h07;
            16'd13858: data <= 8'hE0;
            16'd13859: data <= 8'h07;
            16'd13860: data <= 8'hE0;
            16'd13861: data <= 8'h07;
            16'd13862: data <= 8'hE0;
            16'd13863: data <= 8'h07;
            16'd13864: data <= 8'hE0;
            16'd13865: data <= 8'h07;
            16'd13866: data <= 8'hE0;
            16'd13867: data <= 8'h07;
            16'd13868: data <= 8'hE0;
            16'd13869: data <= 8'h07;
            16'd13870: data <= 8'hE0;
            16'd13871: data <= 8'h07;
            16'd13872: data <= 8'hE0;
            16'd13873: data <= 8'h07;
            16'd13874: data <= 8'hE0;
            16'd13875: data <= 8'h07;
            16'd13876: data <= 8'hE0;
            16'd13877: data <= 8'h07;
            16'd13878: data <= 8'hE0;
            16'd13879: data <= 8'h07;
            16'd13880: data <= 8'hFF;
            16'd13881: data <= 8'hFF;
            16'd13882: data <= 8'hE0;
            16'd13883: data <= 8'h07;
            16'd13884: data <= 8'hE0;
            16'd13885: data <= 8'h07;
            16'd13886: data <= 8'hE0;
            16'd13887: data <= 8'h07;
            16'd13888: data <= 8'hE0;
            16'd13889: data <= 8'h07;
            16'd13890: data <= 8'hE0;
            16'd13891: data <= 8'h07;
            16'd13892: data <= 8'hE0;
            16'd13893: data <= 8'h07;
            16'd13894: data <= 8'hE0;
            16'd13895: data <= 8'h07;
            16'd13896: data <= 8'hE0;
            16'd13897: data <= 8'h07;
            16'd13898: data <= 8'hE0;
            16'd13899: data <= 8'h07;
            16'd13900: data <= 8'hE0;
            16'd13901: data <= 8'h07;
            16'd13902: data <= 8'hE0;
            16'd13903: data <= 8'h07;
            16'd13904: data <= 8'hE0;
            16'd13905: data <= 8'h07;
            16'd13906: data <= 8'hE0;
            16'd13907: data <= 8'h07;
            16'd13908: data <= 8'hE0;
            16'd13909: data <= 8'h07;
            16'd13910: data <= 8'hE0;
            16'd13911: data <= 8'h07;
            16'd13912: data <= 8'hE0;
            16'd13913: data <= 8'h07;
            16'd13914: data <= 8'hE0;
            16'd13915: data <= 8'h07;
            16'd13916: data <= 8'hE0;
            16'd13917: data <= 8'h07;
            16'd13918: data <= 8'hE0;
            16'd13919: data <= 8'h07;
            16'd13920: data <= 8'hFF;
            16'd13921: data <= 8'hFF;
            16'd13922: data <= 8'hE0;
            16'd13923: data <= 8'h07;
            16'd13924: data <= 8'hE0;
            16'd13925: data <= 8'h07;
            16'd13926: data <= 8'hE0;
            16'd13927: data <= 8'h07;
            16'd13928: data <= 8'hE0;
            16'd13929: data <= 8'h07;
            16'd13930: data <= 8'hE0;
            16'd13931: data <= 8'h07;
            16'd13932: data <= 8'hE0;
            16'd13933: data <= 8'h07;
            16'd13934: data <= 8'hE0;
            16'd13935: data <= 8'h07;
            16'd13936: data <= 8'hE0;
            16'd13937: data <= 8'h07;
            16'd13938: data <= 8'hE0;
            16'd13939: data <= 8'h07;
            16'd13940: data <= 8'hE0;
            16'd13941: data <= 8'h07;
            16'd13942: data <= 8'hE0;
            16'd13943: data <= 8'h07;
            16'd13944: data <= 8'hE0;
            16'd13945: data <= 8'h07;
            16'd13946: data <= 8'hE0;
            16'd13947: data <= 8'h07;
            16'd13948: data <= 8'hE0;
            16'd13949: data <= 8'h07;
            16'd13950: data <= 8'hE0;
            16'd13951: data <= 8'h07;
            16'd13952: data <= 8'hE0;
            16'd13953: data <= 8'h07;
            16'd13954: data <= 8'hE0;
            16'd13955: data <= 8'h07;
            16'd13956: data <= 8'hE0;
            16'd13957: data <= 8'h07;
            16'd13958: data <= 8'hE0;
            16'd13959: data <= 8'h07;
            16'd13960: data <= 8'hFF;
            16'd13961: data <= 8'hFF;
            16'd13962: data <= 8'hE0;
            16'd13963: data <= 8'h07;
            16'd13964: data <= 8'hE0;
            16'd13965: data <= 8'h07;
            16'd13966: data <= 8'hE0;
            16'd13967: data <= 8'h07;
            16'd13968: data <= 8'hE0;
            16'd13969: data <= 8'h07;
            16'd13970: data <= 8'hE0;
            16'd13971: data <= 8'h07;
            16'd13972: data <= 8'hE0;
            16'd13973: data <= 8'h07;
            16'd13974: data <= 8'hE0;
            16'd13975: data <= 8'h07;
            16'd13976: data <= 8'hE0;
            16'd13977: data <= 8'h07;
            16'd13978: data <= 8'hE0;
            16'd13979: data <= 8'h07;
            16'd13980: data <= 8'hE0;
            16'd13981: data <= 8'h07;
            16'd13982: data <= 8'hE0;
            16'd13983: data <= 8'h07;
            16'd13984: data <= 8'hE0;
            16'd13985: data <= 8'h07;
            16'd13986: data <= 8'hE0;
            16'd13987: data <= 8'h07;
            16'd13988: data <= 8'hE0;
            16'd13989: data <= 8'h07;
            16'd13990: data <= 8'hE0;
            16'd13991: data <= 8'h07;
            16'd13992: data <= 8'hE0;
            16'd13993: data <= 8'h07;
            16'd13994: data <= 8'hE0;
            16'd13995: data <= 8'h07;
            16'd13996: data <= 8'hE0;
            16'd13997: data <= 8'h07;
            16'd13998: data <= 8'hE0;
            16'd13999: data <= 8'h07;
            16'd14000: data <= 8'hFF;
            16'd14001: data <= 8'hFF;
            16'd14002: data <= 8'hE0;
            16'd14003: data <= 8'h07;
            16'd14004: data <= 8'hE0;
            16'd14005: data <= 8'h07;
            16'd14006: data <= 8'hE0;
            16'd14007: data <= 8'h07;
            16'd14008: data <= 8'hE0;
            16'd14009: data <= 8'h07;
            16'd14010: data <= 8'hE0;
            16'd14011: data <= 8'h07;
            16'd14012: data <= 8'hE0;
            16'd14013: data <= 8'h07;
            16'd14014: data <= 8'hE0;
            16'd14015: data <= 8'h07;
            16'd14016: data <= 8'hE0;
            16'd14017: data <= 8'h07;
            16'd14018: data <= 8'hE0;
            16'd14019: data <= 8'h07;
            16'd14020: data <= 8'hE0;
            16'd14021: data <= 8'h07;
            16'd14022: data <= 8'hE0;
            16'd14023: data <= 8'h07;
            16'd14024: data <= 8'hE0;
            16'd14025: data <= 8'h07;
            16'd14026: data <= 8'hE0;
            16'd14027: data <= 8'h07;
            16'd14028: data <= 8'hE0;
            16'd14029: data <= 8'h07;
            16'd14030: data <= 8'hE0;
            16'd14031: data <= 8'h07;
            16'd14032: data <= 8'hE0;
            16'd14033: data <= 8'h07;
            16'd14034: data <= 8'hE0;
            16'd14035: data <= 8'h07;
            16'd14036: data <= 8'hE0;
            16'd14037: data <= 8'h07;
            16'd14038: data <= 8'hE0;
            16'd14039: data <= 8'h07;
            16'd14040: data <= 8'hFF;
            16'd14041: data <= 8'hFF;
            16'd14042: data <= 8'hE0;
            16'd14043: data <= 8'h07;
            16'd14044: data <= 8'hE0;
            16'd14045: data <= 8'h07;
            16'd14046: data <= 8'hE0;
            16'd14047: data <= 8'h07;
            16'd14048: data <= 8'hE0;
            16'd14049: data <= 8'h07;
            16'd14050: data <= 8'hE0;
            16'd14051: data <= 8'h07;
            16'd14052: data <= 8'hE0;
            16'd14053: data <= 8'h07;
            16'd14054: data <= 8'hE0;
            16'd14055: data <= 8'h07;
            16'd14056: data <= 8'hE0;
            16'd14057: data <= 8'h07;
            16'd14058: data <= 8'hE0;
            16'd14059: data <= 8'h07;
            16'd14060: data <= 8'hE0;
            16'd14061: data <= 8'h07;
            16'd14062: data <= 8'hE0;
            16'd14063: data <= 8'h07;
            16'd14064: data <= 8'hE0;
            16'd14065: data <= 8'h07;
            16'd14066: data <= 8'hE0;
            16'd14067: data <= 8'h07;
            16'd14068: data <= 8'hE0;
            16'd14069: data <= 8'h07;
            16'd14070: data <= 8'hE0;
            16'd14071: data <= 8'h07;
            16'd14072: data <= 8'hE0;
            16'd14073: data <= 8'h07;
            16'd14074: data <= 8'hE0;
            16'd14075: data <= 8'h07;
            16'd14076: data <= 8'hE0;
            16'd14077: data <= 8'h07;
            16'd14078: data <= 8'hE0;
            16'd14079: data <= 8'h07;
            16'd14080: data <= 8'hFF;
            16'd14081: data <= 8'hFF;
            16'd14082: data <= 8'hE0;
            16'd14083: data <= 8'h07;
            16'd14084: data <= 8'hE0;
            16'd14085: data <= 8'h07;
            16'd14086: data <= 8'hE0;
            16'd14087: data <= 8'h07;
            16'd14088: data <= 8'hE0;
            16'd14089: data <= 8'h07;
            16'd14090: data <= 8'hE0;
            16'd14091: data <= 8'h07;
            16'd14092: data <= 8'hE0;
            16'd14093: data <= 8'h07;
            16'd14094: data <= 8'hE0;
            16'd14095: data <= 8'h07;
            16'd14096: data <= 8'hE0;
            16'd14097: data <= 8'h07;
            16'd14098: data <= 8'hE0;
            16'd14099: data <= 8'h07;
            16'd14100: data <= 8'hE0;
            16'd14101: data <= 8'h07;
            16'd14102: data <= 8'hE0;
            16'd14103: data <= 8'h07;
            16'd14104: data <= 8'hE0;
            16'd14105: data <= 8'h07;
            16'd14106: data <= 8'hE0;
            16'd14107: data <= 8'h07;
            16'd14108: data <= 8'hE0;
            16'd14109: data <= 8'h07;
            16'd14110: data <= 8'hE0;
            16'd14111: data <= 8'h07;
            16'd14112: data <= 8'hE0;
            16'd14113: data <= 8'h07;
            16'd14114: data <= 8'hE0;
            16'd14115: data <= 8'h07;
            16'd14116: data <= 8'hE0;
            16'd14117: data <= 8'h07;
            16'd14118: data <= 8'hE0;
            16'd14119: data <= 8'h07;
            16'd14120: data <= 8'hFF;
            16'd14121: data <= 8'hFF;
            16'd14122: data <= 8'hE0;
            16'd14123: data <= 8'h07;
            16'd14124: data <= 8'hE0;
            16'd14125: data <= 8'h07;
            16'd14126: data <= 8'hE0;
            16'd14127: data <= 8'h07;
            16'd14128: data <= 8'hE0;
            16'd14129: data <= 8'h07;
            16'd14130: data <= 8'hE0;
            16'd14131: data <= 8'h07;
            16'd14132: data <= 8'hE0;
            16'd14133: data <= 8'h07;
            16'd14134: data <= 8'hE0;
            16'd14135: data <= 8'h07;
            16'd14136: data <= 8'hE0;
            16'd14137: data <= 8'h07;
            16'd14138: data <= 8'hE0;
            16'd14139: data <= 8'h07;
            16'd14140: data <= 8'hE0;
            16'd14141: data <= 8'h07;
            16'd14142: data <= 8'hE0;
            16'd14143: data <= 8'h07;
            16'd14144: data <= 8'hE0;
            16'd14145: data <= 8'h07;
            16'd14146: data <= 8'hE0;
            16'd14147: data <= 8'h07;
            16'd14148: data <= 8'hE0;
            16'd14149: data <= 8'h07;
            16'd14150: data <= 8'hE0;
            16'd14151: data <= 8'h07;
            16'd14152: data <= 8'hE0;
            16'd14153: data <= 8'h07;
            16'd14154: data <= 8'hE0;
            16'd14155: data <= 8'h07;
            16'd14156: data <= 8'hE0;
            16'd14157: data <= 8'h07;
            16'd14158: data <= 8'hE0;
            16'd14159: data <= 8'h07;
            16'd14160: data <= 8'hFF;
            16'd14161: data <= 8'hFF;
            16'd14162: data <= 8'hE0;
            16'd14163: data <= 8'h07;
            16'd14164: data <= 8'hE0;
            16'd14165: data <= 8'h07;
            16'd14166: data <= 8'hE0;
            16'd14167: data <= 8'h07;
            16'd14168: data <= 8'hE0;
            16'd14169: data <= 8'h07;
            16'd14170: data <= 8'hE0;
            16'd14171: data <= 8'h07;
            16'd14172: data <= 8'hE0;
            16'd14173: data <= 8'h07;
            16'd14174: data <= 8'hE0;
            16'd14175: data <= 8'h07;
            16'd14176: data <= 8'hE0;
            16'd14177: data <= 8'h07;
            16'd14178: data <= 8'hE0;
            16'd14179: data <= 8'h07;
            16'd14180: data <= 8'hE0;
            16'd14181: data <= 8'h07;
            16'd14182: data <= 8'hE0;
            16'd14183: data <= 8'h07;
            16'd14184: data <= 8'hE0;
            16'd14185: data <= 8'h07;
            16'd14186: data <= 8'hE0;
            16'd14187: data <= 8'h07;
            16'd14188: data <= 8'hE0;
            16'd14189: data <= 8'h07;
            16'd14190: data <= 8'hE0;
            16'd14191: data <= 8'h07;
            16'd14192: data <= 8'hE0;
            16'd14193: data <= 8'h07;
            16'd14194: data <= 8'hE0;
            16'd14195: data <= 8'h07;
            16'd14196: data <= 8'hE0;
            16'd14197: data <= 8'h07;
            16'd14198: data <= 8'hE0;
            16'd14199: data <= 8'h07;
            16'd14200: data <= 8'hFF;
            16'd14201: data <= 8'hFF;
            16'd14202: data <= 8'hE0;
            16'd14203: data <= 8'h07;
            16'd14204: data <= 8'hE0;
            16'd14205: data <= 8'h07;
            16'd14206: data <= 8'hE0;
            16'd14207: data <= 8'h07;
            16'd14208: data <= 8'hE0;
            16'd14209: data <= 8'h07;
            16'd14210: data <= 8'hE0;
            16'd14211: data <= 8'h07;
            16'd14212: data <= 8'hE0;
            16'd14213: data <= 8'h07;
            16'd14214: data <= 8'hE0;
            16'd14215: data <= 8'h07;
            16'd14216: data <= 8'hE0;
            16'd14217: data <= 8'h07;
            16'd14218: data <= 8'hE0;
            16'd14219: data <= 8'h07;
            16'd14220: data <= 8'hE0;
            16'd14221: data <= 8'h07;
            16'd14222: data <= 8'hE0;
            16'd14223: data <= 8'h07;
            16'd14224: data <= 8'hE0;
            16'd14225: data <= 8'h07;
            16'd14226: data <= 8'hE0;
            16'd14227: data <= 8'h07;
            16'd14228: data <= 8'hE0;
            16'd14229: data <= 8'h07;
            16'd14230: data <= 8'hE0;
            16'd14231: data <= 8'h07;
            16'd14232: data <= 8'hE0;
            16'd14233: data <= 8'h07;
            16'd14234: data <= 8'hE0;
            16'd14235: data <= 8'h07;
            16'd14236: data <= 8'hE0;
            16'd14237: data <= 8'h07;
            16'd14238: data <= 8'hE0;
            16'd14239: data <= 8'h07;
            16'd14240: data <= 8'hFF;
            16'd14241: data <= 8'hFF;
            16'd14242: data <= 8'hE0;
            16'd14243: data <= 8'h07;
            16'd14244: data <= 8'hE0;
            16'd14245: data <= 8'h07;
            16'd14246: data <= 8'hE0;
            16'd14247: data <= 8'h07;
            16'd14248: data <= 8'hE0;
            16'd14249: data <= 8'h07;
            16'd14250: data <= 8'hE0;
            16'd14251: data <= 8'h07;
            16'd14252: data <= 8'hE0;
            16'd14253: data <= 8'h07;
            16'd14254: data <= 8'hE0;
            16'd14255: data <= 8'h07;
            16'd14256: data <= 8'hE0;
            16'd14257: data <= 8'h07;
            16'd14258: data <= 8'hE0;
            16'd14259: data <= 8'h07;
            16'd14260: data <= 8'hE0;
            16'd14261: data <= 8'h07;
            16'd14262: data <= 8'hE0;
            16'd14263: data <= 8'h07;
            16'd14264: data <= 8'hE0;
            16'd14265: data <= 8'h07;
            16'd14266: data <= 8'hE0;
            16'd14267: data <= 8'h07;
            16'd14268: data <= 8'hE0;
            16'd14269: data <= 8'h07;
            16'd14270: data <= 8'hE0;
            16'd14271: data <= 8'h07;
            16'd14272: data <= 8'hE0;
            16'd14273: data <= 8'h07;
            16'd14274: data <= 8'hE0;
            16'd14275: data <= 8'h07;
            16'd14276: data <= 8'hE0;
            16'd14277: data <= 8'h07;
            16'd14278: data <= 8'hE0;
            16'd14279: data <= 8'h07;
            16'd14280: data <= 8'hFF;
            16'd14281: data <= 8'hFF;
            16'd14282: data <= 8'hE0;
            16'd14283: data <= 8'h07;
            16'd14284: data <= 8'hE0;
            16'd14285: data <= 8'h07;
            16'd14286: data <= 8'hE0;
            16'd14287: data <= 8'h07;
            16'd14288: data <= 8'hE0;
            16'd14289: data <= 8'h07;
            16'd14290: data <= 8'hE0;
            16'd14291: data <= 8'h07;
            16'd14292: data <= 8'hE0;
            16'd14293: data <= 8'h07;
            16'd14294: data <= 8'hE0;
            16'd14295: data <= 8'h07;
            16'd14296: data <= 8'hE0;
            16'd14297: data <= 8'h07;
            16'd14298: data <= 8'hE0;
            16'd14299: data <= 8'h07;
            16'd14300: data <= 8'hE0;
            16'd14301: data <= 8'h07;
            16'd14302: data <= 8'hE0;
            16'd14303: data <= 8'h07;
            16'd14304: data <= 8'hE0;
            16'd14305: data <= 8'h07;
            16'd14306: data <= 8'hE0;
            16'd14307: data <= 8'h07;
            16'd14308: data <= 8'hE0;
            16'd14309: data <= 8'h07;
            16'd14310: data <= 8'hE0;
            16'd14311: data <= 8'h07;
            16'd14312: data <= 8'hE0;
            16'd14313: data <= 8'h07;
            16'd14314: data <= 8'hE0;
            16'd14315: data <= 8'h07;
            16'd14316: data <= 8'hE0;
            16'd14317: data <= 8'h07;
            16'd14318: data <= 8'hE0;
            16'd14319: data <= 8'h07;
            16'd14320: data <= 8'hFF;
            16'd14321: data <= 8'hFF;
            16'd14322: data <= 8'hE0;
            16'd14323: data <= 8'h07;
            16'd14324: data <= 8'hE0;
            16'd14325: data <= 8'h07;
            16'd14326: data <= 8'hE0;
            16'd14327: data <= 8'h07;
            16'd14328: data <= 8'hE0;
            16'd14329: data <= 8'h07;
            16'd14330: data <= 8'hE0;
            16'd14331: data <= 8'h07;
            16'd14332: data <= 8'hE0;
            16'd14333: data <= 8'h07;
            16'd14334: data <= 8'hE0;
            16'd14335: data <= 8'h07;
            16'd14336: data <= 8'hE0;
            16'd14337: data <= 8'h07;
            16'd14338: data <= 8'hE0;
            16'd14339: data <= 8'h07;
            16'd14340: data <= 8'hE0;
            16'd14341: data <= 8'h07;
            16'd14342: data <= 8'hE0;
            16'd14343: data <= 8'h07;
            16'd14344: data <= 8'hE0;
            16'd14345: data <= 8'h07;
            16'd14346: data <= 8'hE0;
            16'd14347: data <= 8'h07;
            16'd14348: data <= 8'hE0;
            16'd14349: data <= 8'h07;
            16'd14350: data <= 8'hE0;
            16'd14351: data <= 8'h07;
            16'd14352: data <= 8'hE0;
            16'd14353: data <= 8'h07;
            16'd14354: data <= 8'hE0;
            16'd14355: data <= 8'h07;
            16'd14356: data <= 8'hE0;
            16'd14357: data <= 8'h07;
            16'd14358: data <= 8'hE0;
            16'd14359: data <= 8'h07;
            16'd14360: data <= 8'hFF;
            16'd14361: data <= 8'hFF;
            16'd14362: data <= 8'hE0;
            16'd14363: data <= 8'h07;
            16'd14364: data <= 8'hE0;
            16'd14365: data <= 8'h07;
            16'd14366: data <= 8'hE0;
            16'd14367: data <= 8'h07;
            16'd14368: data <= 8'hE0;
            16'd14369: data <= 8'h07;
            16'd14370: data <= 8'hE0;
            16'd14371: data <= 8'h07;
            16'd14372: data <= 8'hE0;
            16'd14373: data <= 8'h07;
            16'd14374: data <= 8'hE0;
            16'd14375: data <= 8'h07;
            16'd14376: data <= 8'hE0;
            16'd14377: data <= 8'h07;
            16'd14378: data <= 8'hE0;
            16'd14379: data <= 8'h07;
            16'd14380: data <= 8'hE0;
            16'd14381: data <= 8'h07;
            16'd14382: data <= 8'hE0;
            16'd14383: data <= 8'h07;
            16'd14384: data <= 8'hE0;
            16'd14385: data <= 8'h07;
            16'd14386: data <= 8'hE0;
            16'd14387: data <= 8'h07;
            16'd14388: data <= 8'hE0;
            16'd14389: data <= 8'h07;
            16'd14390: data <= 8'hE0;
            16'd14391: data <= 8'h07;
            16'd14392: data <= 8'hE0;
            16'd14393: data <= 8'h07;
            16'd14394: data <= 8'hE0;
            16'd14395: data <= 8'h07;
            16'd14396: data <= 8'hE0;
            16'd14397: data <= 8'h07;
            16'd14398: data <= 8'hE0;
            16'd14399: data <= 8'h07;
            16'd14400: data <= 8'hFF;
            16'd14401: data <= 8'hFF;
            16'd14402: data <= 8'hFF;
            16'd14403: data <= 8'hFF;
            16'd14404: data <= 8'hFF;
            16'd14405: data <= 8'hFF;
            16'd14406: data <= 8'hFF;
            16'd14407: data <= 8'hFF;
            16'd14408: data <= 8'hFF;
            16'd14409: data <= 8'hFF;
            16'd14410: data <= 8'hFF;
            16'd14411: data <= 8'hFF;
            16'd14412: data <= 8'hFF;
            16'd14413: data <= 8'hFF;
            16'd14414: data <= 8'hFF;
            16'd14415: data <= 8'hFF;
            16'd14416: data <= 8'hFF;
            16'd14417: data <= 8'hFF;
            16'd14418: data <= 8'hFF;
            16'd14419: data <= 8'hFF;
            16'd14420: data <= 8'hFF;
            16'd14421: data <= 8'hFF;
            16'd14422: data <= 8'hFF;
            16'd14423: data <= 8'hFF;
            16'd14424: data <= 8'hFF;
            16'd14425: data <= 8'hFF;
            16'd14426: data <= 8'hFF;
            16'd14427: data <= 8'hFF;
            16'd14428: data <= 8'hFF;
            16'd14429: data <= 8'hFF;
            16'd14430: data <= 8'hFF;
            16'd14431: data <= 8'hFF;
            16'd14432: data <= 8'hFF;
            16'd14433: data <= 8'hFF;
            16'd14434: data <= 8'hFF;
            16'd14435: data <= 8'hFF;
            16'd14436: data <= 8'hFF;
            16'd14437: data <= 8'hFF;
            16'd14438: data <= 8'hFF;
            16'd14439: data <= 8'hFF;
            16'd14440: data <= 8'hFF;
            16'd14441: data <= 8'hFF;
            16'd14442: data <= 8'hFF;
            16'd14443: data <= 8'hFF;
            16'd14444: data <= 8'hFF;
            16'd14445: data <= 8'hFF;
            16'd14446: data <= 8'hFF;
            16'd14447: data <= 8'hFF;
            16'd14448: data <= 8'hFF;
            16'd14449: data <= 8'hFF;
            16'd14450: data <= 8'hFF;
            16'd14451: data <= 8'hFF;
            16'd14452: data <= 8'hFF;
            16'd14453: data <= 8'hFF;
            16'd14454: data <= 8'hFF;
            16'd14455: data <= 8'hFF;
            16'd14456: data <= 8'hFF;
            16'd14457: data <= 8'hFF;
            16'd14458: data <= 8'hFF;
            16'd14459: data <= 8'hFF;
            16'd14460: data <= 8'hFF;
            16'd14461: data <= 8'hFF;
            16'd14462: data <= 8'hFF;
            16'd14463: data <= 8'hFF;
            16'd14464: data <= 8'hFF;
            16'd14465: data <= 8'hFF;
            16'd14466: data <= 8'hFF;
            16'd14467: data <= 8'hFF;
            16'd14468: data <= 8'hFF;
            16'd14469: data <= 8'hFF;
            16'd14470: data <= 8'hFF;
            16'd14471: data <= 8'hFF;
            16'd14472: data <= 8'hFF;
            16'd14473: data <= 8'hFF;
            16'd14474: data <= 8'hFF;
            16'd14475: data <= 8'hFF;
            16'd14476: data <= 8'hFF;
            16'd14477: data <= 8'hFF;
            16'd14478: data <= 8'hFF;
            16'd14479: data <= 8'hFF;
            16'd14480: data <= 8'hFF;
            16'd14481: data <= 8'hFF;
            16'd14482: data <= 8'hFF;
            16'd14483: data <= 8'hFF;
            16'd14484: data <= 8'hFF;
            16'd14485: data <= 8'hFF;
            16'd14486: data <= 8'hFF;
            16'd14487: data <= 8'hFF;
            16'd14488: data <= 8'hFF;
            16'd14489: data <= 8'hFF;
            16'd14490: data <= 8'hFF;
            16'd14491: data <= 8'hFF;
            16'd14492: data <= 8'hFF;
            16'd14493: data <= 8'hFF;
            16'd14494: data <= 8'hFF;
            16'd14495: data <= 8'hFF;
            16'd14496: data <= 8'hFF;
            16'd14497: data <= 8'hFF;
            16'd14498: data <= 8'hFF;
            16'd14499: data <= 8'hFF;
            16'd14500: data <= 8'hFF;
            16'd14501: data <= 8'hFF;
            16'd14502: data <= 8'hFF;
            16'd14503: data <= 8'hFF;
            16'd14504: data <= 8'hFF;
            16'd14505: data <= 8'hFF;
            16'd14506: data <= 8'hFF;
            16'd14507: data <= 8'hFF;
            16'd14508: data <= 8'hFF;
            16'd14509: data <= 8'hFF;
            16'd14510: data <= 8'hFF;
            16'd14511: data <= 8'hFF;
            16'd14512: data <= 8'hFF;
            16'd14513: data <= 8'hFF;
            16'd14514: data <= 8'hFF;
            16'd14515: data <= 8'hFF;
            16'd14516: data <= 8'hFF;
            16'd14517: data <= 8'hFF;
            16'd14518: data <= 8'hFF;
            16'd14519: data <= 8'hFF;
            16'd14520: data <= 8'hFF;
            16'd14521: data <= 8'hFF;
            16'd14522: data <= 8'hFF;
            16'd14523: data <= 8'hFF;
            16'd14524: data <= 8'hFF;
            16'd14525: data <= 8'hFF;
            16'd14526: data <= 8'hFF;
            16'd14527: data <= 8'hFF;
            16'd14528: data <= 8'hFF;
            16'd14529: data <= 8'hFF;
            16'd14530: data <= 8'hFF;
            16'd14531: data <= 8'hFF;
            16'd14532: data <= 8'hFF;
            16'd14533: data <= 8'hFF;
            16'd14534: data <= 8'hFF;
            16'd14535: data <= 8'hFF;
            16'd14536: data <= 8'hFF;
            16'd14537: data <= 8'hFF;
            16'd14538: data <= 8'hFF;
            16'd14539: data <= 8'hFF;
            16'd14540: data <= 8'hFF;
            16'd14541: data <= 8'hFF;
            16'd14542: data <= 8'hFF;
            16'd14543: data <= 8'hFF;
            16'd14544: data <= 8'hFF;
            16'd14545: data <= 8'hFF;
            16'd14546: data <= 8'hFF;
            16'd14547: data <= 8'hFF;
            16'd14548: data <= 8'hFF;
            16'd14549: data <= 8'hFF;
            16'd14550: data <= 8'hFF;
            16'd14551: data <= 8'hFF;
            16'd14552: data <= 8'hFF;
            16'd14553: data <= 8'hFF;
            16'd14554: data <= 8'hFF;
            16'd14555: data <= 8'hFF;
            16'd14556: data <= 8'hFF;
            16'd14557: data <= 8'hFF;
            16'd14558: data <= 8'hFF;
            16'd14559: data <= 8'hFF;
            16'd14560: data <= 8'hFF;
            16'd14561: data <= 8'hFF;
            16'd14562: data <= 8'hFF;
            16'd14563: data <= 8'hFF;
            16'd14564: data <= 8'hFF;
            16'd14565: data <= 8'hFF;
            16'd14566: data <= 8'hFF;
            16'd14567: data <= 8'hFF;
            16'd14568: data <= 8'hFF;
            16'd14569: data <= 8'hFF;
            16'd14570: data <= 8'hFF;
            16'd14571: data <= 8'hFF;
            16'd14572: data <= 8'hFF;
            16'd14573: data <= 8'hFF;
            16'd14574: data <= 8'hFF;
            16'd14575: data <= 8'hFF;
            16'd14576: data <= 8'hFF;
            16'd14577: data <= 8'hFF;
            16'd14578: data <= 8'hFF;
            16'd14579: data <= 8'hFF;
            16'd14580: data <= 8'hFF;
            16'd14581: data <= 8'hFF;
            16'd14582: data <= 8'hFF;
            16'd14583: data <= 8'hFF;
            16'd14584: data <= 8'hFF;
            16'd14585: data <= 8'hFF;
            16'd14586: data <= 8'hFF;
            16'd14587: data <= 8'hFF;
            16'd14588: data <= 8'hFF;
            16'd14589: data <= 8'hFF;
            16'd14590: data <= 8'hFF;
            16'd14591: data <= 8'hFF;
            16'd14592: data <= 8'hFF;
            16'd14593: data <= 8'hFF;
            16'd14594: data <= 8'hFF;
            16'd14595: data <= 8'hFF;
            16'd14596: data <= 8'hFF;
            16'd14597: data <= 8'hFF;
            16'd14598: data <= 8'hFF;
            16'd14599: data <= 8'hFF;
            16'd14600: data <= 8'hFF;
            16'd14601: data <= 8'hFF;
            16'd14602: data <= 8'hFF;
            16'd14603: data <= 8'hFF;
            16'd14604: data <= 8'hFF;
            16'd14605: data <= 8'hFF;
            16'd14606: data <= 8'hFF;
            16'd14607: data <= 8'hFF;
            16'd14608: data <= 8'hFF;
            16'd14609: data <= 8'hFF;
            16'd14610: data <= 8'hFF;
            16'd14611: data <= 8'hFF;
            16'd14612: data <= 8'hFF;
            16'd14613: data <= 8'hFF;
            16'd14614: data <= 8'hFF;
            16'd14615: data <= 8'hFF;
            16'd14616: data <= 8'hFF;
            16'd14617: data <= 8'hFF;
            16'd14618: data <= 8'hFF;
            16'd14619: data <= 8'hFF;
            16'd14620: data <= 8'hFF;
            16'd14621: data <= 8'hFF;
            16'd14622: data <= 8'hFF;
            16'd14623: data <= 8'hFF;
            16'd14624: data <= 8'hFF;
            16'd14625: data <= 8'hFF;
            16'd14626: data <= 8'hFF;
            16'd14627: data <= 8'hFF;
            16'd14628: data <= 8'hFF;
            16'd14629: data <= 8'hFF;
            16'd14630: data <= 8'hFF;
            16'd14631: data <= 8'hFF;
            16'd14632: data <= 8'hFF;
            16'd14633: data <= 8'hFF;
            16'd14634: data <= 8'hFF;
            16'd14635: data <= 8'hFF;
            16'd14636: data <= 8'hFF;
            16'd14637: data <= 8'hFF;
            16'd14638: data <= 8'hFF;
            16'd14639: data <= 8'hFF;
            16'd14640: data <= 8'hFF;
            16'd14641: data <= 8'hFF;
            16'd14642: data <= 8'hE0;
            16'd14643: data <= 8'h07;
            16'd14644: data <= 8'hE0;
            16'd14645: data <= 8'h07;
            16'd14646: data <= 8'hE0;
            16'd14647: data <= 8'h07;
            16'd14648: data <= 8'hE0;
            16'd14649: data <= 8'h07;
            16'd14650: data <= 8'hE0;
            16'd14651: data <= 8'h07;
            16'd14652: data <= 8'hE0;
            16'd14653: data <= 8'h07;
            16'd14654: data <= 8'hE0;
            16'd14655: data <= 8'h07;
            16'd14656: data <= 8'hE0;
            16'd14657: data <= 8'h07;
            16'd14658: data <= 8'hE0;
            16'd14659: data <= 8'h07;
            16'd14660: data <= 8'hE0;
            16'd14661: data <= 8'h07;
            16'd14662: data <= 8'hE0;
            16'd14663: data <= 8'h07;
            16'd14664: data <= 8'hE0;
            16'd14665: data <= 8'h07;
            16'd14666: data <= 8'hE0;
            16'd14667: data <= 8'h07;
            16'd14668: data <= 8'hE0;
            16'd14669: data <= 8'h07;
            16'd14670: data <= 8'hE0;
            16'd14671: data <= 8'h07;
            16'd14672: data <= 8'hE0;
            16'd14673: data <= 8'h07;
            16'd14674: data <= 8'hE0;
            16'd14675: data <= 8'h07;
            16'd14676: data <= 8'hE0;
            16'd14677: data <= 8'h07;
            16'd14678: data <= 8'hE0;
            16'd14679: data <= 8'h07;
            16'd14680: data <= 8'hFF;
            16'd14681: data <= 8'hFF;
            16'd14682: data <= 8'hE0;
            16'd14683: data <= 8'h07;
            16'd14684: data <= 8'hE0;
            16'd14685: data <= 8'h07;
            16'd14686: data <= 8'hE0;
            16'd14687: data <= 8'h07;
            16'd14688: data <= 8'hE0;
            16'd14689: data <= 8'h07;
            16'd14690: data <= 8'hE0;
            16'd14691: data <= 8'h07;
            16'd14692: data <= 8'hE0;
            16'd14693: data <= 8'h07;
            16'd14694: data <= 8'hE0;
            16'd14695: data <= 8'h07;
            16'd14696: data <= 8'hE0;
            16'd14697: data <= 8'h07;
            16'd14698: data <= 8'hE0;
            16'd14699: data <= 8'h07;
            16'd14700: data <= 8'hE0;
            16'd14701: data <= 8'h07;
            16'd14702: data <= 8'hE0;
            16'd14703: data <= 8'h07;
            16'd14704: data <= 8'hE0;
            16'd14705: data <= 8'h07;
            16'd14706: data <= 8'hE0;
            16'd14707: data <= 8'h07;
            16'd14708: data <= 8'hE0;
            16'd14709: data <= 8'h07;
            16'd14710: data <= 8'hE0;
            16'd14711: data <= 8'h07;
            16'd14712: data <= 8'hE0;
            16'd14713: data <= 8'h07;
            16'd14714: data <= 8'hE0;
            16'd14715: data <= 8'h07;
            16'd14716: data <= 8'hE0;
            16'd14717: data <= 8'h07;
            16'd14718: data <= 8'hE0;
            16'd14719: data <= 8'h07;
            16'd14720: data <= 8'hFF;
            16'd14721: data <= 8'hFF;
            16'd14722: data <= 8'hE0;
            16'd14723: data <= 8'h07;
            16'd14724: data <= 8'hE0;
            16'd14725: data <= 8'h07;
            16'd14726: data <= 8'hE0;
            16'd14727: data <= 8'h07;
            16'd14728: data <= 8'hE0;
            16'd14729: data <= 8'h07;
            16'd14730: data <= 8'hE0;
            16'd14731: data <= 8'h07;
            16'd14732: data <= 8'hE0;
            16'd14733: data <= 8'h07;
            16'd14734: data <= 8'hE0;
            16'd14735: data <= 8'h07;
            16'd14736: data <= 8'hE0;
            16'd14737: data <= 8'h07;
            16'd14738: data <= 8'hE0;
            16'd14739: data <= 8'h07;
            16'd14740: data <= 8'hE0;
            16'd14741: data <= 8'h07;
            16'd14742: data <= 8'hE0;
            16'd14743: data <= 8'h07;
            16'd14744: data <= 8'hE0;
            16'd14745: data <= 8'h07;
            16'd14746: data <= 8'hE0;
            16'd14747: data <= 8'h07;
            16'd14748: data <= 8'hE0;
            16'd14749: data <= 8'h07;
            16'd14750: data <= 8'hE0;
            16'd14751: data <= 8'h07;
            16'd14752: data <= 8'hE0;
            16'd14753: data <= 8'h07;
            16'd14754: data <= 8'hE0;
            16'd14755: data <= 8'h07;
            16'd14756: data <= 8'hE0;
            16'd14757: data <= 8'h07;
            16'd14758: data <= 8'hE0;
            16'd14759: data <= 8'h07;
            16'd14760: data <= 8'hFF;
            16'd14761: data <= 8'hFF;
            16'd14762: data <= 8'hE0;
            16'd14763: data <= 8'h07;
            16'd14764: data <= 8'hE0;
            16'd14765: data <= 8'h07;
            16'd14766: data <= 8'hE0;
            16'd14767: data <= 8'h07;
            16'd14768: data <= 8'hE0;
            16'd14769: data <= 8'h07;
            16'd14770: data <= 8'hE0;
            16'd14771: data <= 8'h07;
            16'd14772: data <= 8'hE0;
            16'd14773: data <= 8'h07;
            16'd14774: data <= 8'hE0;
            16'd14775: data <= 8'h07;
            16'd14776: data <= 8'hE0;
            16'd14777: data <= 8'h07;
            16'd14778: data <= 8'hE0;
            16'd14779: data <= 8'h07;
            16'd14780: data <= 8'hE0;
            16'd14781: data <= 8'h07;
            16'd14782: data <= 8'hE0;
            16'd14783: data <= 8'h07;
            16'd14784: data <= 8'hE0;
            16'd14785: data <= 8'h07;
            16'd14786: data <= 8'hE0;
            16'd14787: data <= 8'h07;
            16'd14788: data <= 8'hE0;
            16'd14789: data <= 8'h07;
            16'd14790: data <= 8'hE0;
            16'd14791: data <= 8'h07;
            16'd14792: data <= 8'hE0;
            16'd14793: data <= 8'h07;
            16'd14794: data <= 8'hE0;
            16'd14795: data <= 8'h07;
            16'd14796: data <= 8'hE0;
            16'd14797: data <= 8'h07;
            16'd14798: data <= 8'hE0;
            16'd14799: data <= 8'h07;
            16'd14800: data <= 8'hFF;
            16'd14801: data <= 8'hFF;
            16'd14802: data <= 8'hE0;
            16'd14803: data <= 8'h07;
            16'd14804: data <= 8'hE0;
            16'd14805: data <= 8'h07;
            16'd14806: data <= 8'hE0;
            16'd14807: data <= 8'h07;
            16'd14808: data <= 8'hE0;
            16'd14809: data <= 8'h07;
            16'd14810: data <= 8'hE0;
            16'd14811: data <= 8'h07;
            16'd14812: data <= 8'hE0;
            16'd14813: data <= 8'h07;
            16'd14814: data <= 8'hE0;
            16'd14815: data <= 8'h07;
            16'd14816: data <= 8'hE0;
            16'd14817: data <= 8'h07;
            16'd14818: data <= 8'hE0;
            16'd14819: data <= 8'h07;
            16'd14820: data <= 8'hE0;
            16'd14821: data <= 8'h07;
            16'd14822: data <= 8'hE0;
            16'd14823: data <= 8'h07;
            16'd14824: data <= 8'hE0;
            16'd14825: data <= 8'h07;
            16'd14826: data <= 8'hE0;
            16'd14827: data <= 8'h07;
            16'd14828: data <= 8'hE0;
            16'd14829: data <= 8'h07;
            16'd14830: data <= 8'hE0;
            16'd14831: data <= 8'h07;
            16'd14832: data <= 8'hE0;
            16'd14833: data <= 8'h07;
            16'd14834: data <= 8'hE0;
            16'd14835: data <= 8'h07;
            16'd14836: data <= 8'hE0;
            16'd14837: data <= 8'h07;
            16'd14838: data <= 8'hE0;
            16'd14839: data <= 8'h07;
            16'd14840: data <= 8'hFF;
            16'd14841: data <= 8'hFF;
            16'd14842: data <= 8'hE0;
            16'd14843: data <= 8'h07;
            16'd14844: data <= 8'hE0;
            16'd14845: data <= 8'h07;
            16'd14846: data <= 8'hE0;
            16'd14847: data <= 8'h07;
            16'd14848: data <= 8'hE0;
            16'd14849: data <= 8'h07;
            16'd14850: data <= 8'hE0;
            16'd14851: data <= 8'h07;
            16'd14852: data <= 8'hE0;
            16'd14853: data <= 8'h07;
            16'd14854: data <= 8'hE0;
            16'd14855: data <= 8'h07;
            16'd14856: data <= 8'hE0;
            16'd14857: data <= 8'h07;
            16'd14858: data <= 8'hE0;
            16'd14859: data <= 8'h07;
            16'd14860: data <= 8'hE0;
            16'd14861: data <= 8'h07;
            16'd14862: data <= 8'hE0;
            16'd14863: data <= 8'h07;
            16'd14864: data <= 8'hE0;
            16'd14865: data <= 8'h07;
            16'd14866: data <= 8'hE0;
            16'd14867: data <= 8'h07;
            16'd14868: data <= 8'hE0;
            16'd14869: data <= 8'h07;
            16'd14870: data <= 8'hE0;
            16'd14871: data <= 8'h07;
            16'd14872: data <= 8'hE0;
            16'd14873: data <= 8'h07;
            16'd14874: data <= 8'hE0;
            16'd14875: data <= 8'h07;
            16'd14876: data <= 8'hE0;
            16'd14877: data <= 8'h07;
            16'd14878: data <= 8'hE0;
            16'd14879: data <= 8'h07;
            16'd14880: data <= 8'hFF;
            16'd14881: data <= 8'hFF;
            16'd14882: data <= 8'hE0;
            16'd14883: data <= 8'h07;
            16'd14884: data <= 8'hE0;
            16'd14885: data <= 8'h07;
            16'd14886: data <= 8'hE0;
            16'd14887: data <= 8'h07;
            16'd14888: data <= 8'hE0;
            16'd14889: data <= 8'h07;
            16'd14890: data <= 8'hE0;
            16'd14891: data <= 8'h07;
            16'd14892: data <= 8'hE0;
            16'd14893: data <= 8'h07;
            16'd14894: data <= 8'hE0;
            16'd14895: data <= 8'h07;
            16'd14896: data <= 8'hE0;
            16'd14897: data <= 8'h07;
            16'd14898: data <= 8'hE0;
            16'd14899: data <= 8'h07;
            16'd14900: data <= 8'hE0;
            16'd14901: data <= 8'h07;
            16'd14902: data <= 8'hE0;
            16'd14903: data <= 8'h07;
            16'd14904: data <= 8'hE0;
            16'd14905: data <= 8'h07;
            16'd14906: data <= 8'hE0;
            16'd14907: data <= 8'h07;
            16'd14908: data <= 8'hE0;
            16'd14909: data <= 8'h07;
            16'd14910: data <= 8'hE0;
            16'd14911: data <= 8'h07;
            16'd14912: data <= 8'hE0;
            16'd14913: data <= 8'h07;
            16'd14914: data <= 8'hE0;
            16'd14915: data <= 8'h07;
            16'd14916: data <= 8'hE0;
            16'd14917: data <= 8'h07;
            16'd14918: data <= 8'hE0;
            16'd14919: data <= 8'h07;
            16'd14920: data <= 8'hFF;
            16'd14921: data <= 8'hFF;
            16'd14922: data <= 8'hE0;
            16'd14923: data <= 8'h07;
            16'd14924: data <= 8'hE0;
            16'd14925: data <= 8'h07;
            16'd14926: data <= 8'hE0;
            16'd14927: data <= 8'h07;
            16'd14928: data <= 8'hE0;
            16'd14929: data <= 8'h07;
            16'd14930: data <= 8'hE0;
            16'd14931: data <= 8'h07;
            16'd14932: data <= 8'hE0;
            16'd14933: data <= 8'h07;
            16'd14934: data <= 8'hE0;
            16'd14935: data <= 8'h07;
            16'd14936: data <= 8'hE0;
            16'd14937: data <= 8'h07;
            16'd14938: data <= 8'hE0;
            16'd14939: data <= 8'h07;
            16'd14940: data <= 8'hE0;
            16'd14941: data <= 8'h07;
            16'd14942: data <= 8'hE0;
            16'd14943: data <= 8'h07;
            16'd14944: data <= 8'hE0;
            16'd14945: data <= 8'h07;
            16'd14946: data <= 8'hE0;
            16'd14947: data <= 8'h07;
            16'd14948: data <= 8'hE0;
            16'd14949: data <= 8'h07;
            16'd14950: data <= 8'hE0;
            16'd14951: data <= 8'h07;
            16'd14952: data <= 8'hE0;
            16'd14953: data <= 8'h07;
            16'd14954: data <= 8'hE0;
            16'd14955: data <= 8'h07;
            16'd14956: data <= 8'hE0;
            16'd14957: data <= 8'h07;
            16'd14958: data <= 8'hE0;
            16'd14959: data <= 8'h07;
            16'd14960: data <= 8'hFF;
            16'd14961: data <= 8'hFF;
            16'd14962: data <= 8'hE0;
            16'd14963: data <= 8'h07;
            16'd14964: data <= 8'hE0;
            16'd14965: data <= 8'h07;
            16'd14966: data <= 8'hE0;
            16'd14967: data <= 8'h07;
            16'd14968: data <= 8'hE0;
            16'd14969: data <= 8'h07;
            16'd14970: data <= 8'hE0;
            16'd14971: data <= 8'h07;
            16'd14972: data <= 8'hE0;
            16'd14973: data <= 8'h07;
            16'd14974: data <= 8'hE0;
            16'd14975: data <= 8'h07;
            16'd14976: data <= 8'hE0;
            16'd14977: data <= 8'h07;
            16'd14978: data <= 8'hE0;
            16'd14979: data <= 8'h07;
            16'd14980: data <= 8'hE0;
            16'd14981: data <= 8'h07;
            16'd14982: data <= 8'hE0;
            16'd14983: data <= 8'h07;
            16'd14984: data <= 8'hE0;
            16'd14985: data <= 8'h07;
            16'd14986: data <= 8'hE0;
            16'd14987: data <= 8'h07;
            16'd14988: data <= 8'hE0;
            16'd14989: data <= 8'h07;
            16'd14990: data <= 8'hE0;
            16'd14991: data <= 8'h07;
            16'd14992: data <= 8'hE0;
            16'd14993: data <= 8'h07;
            16'd14994: data <= 8'hE0;
            16'd14995: data <= 8'h07;
            16'd14996: data <= 8'hE0;
            16'd14997: data <= 8'h07;
            16'd14998: data <= 8'hE0;
            16'd14999: data <= 8'h07;
            16'd15000: data <= 8'hFF;
            16'd15001: data <= 8'hFF;
            16'd15002: data <= 8'hE0;
            16'd15003: data <= 8'h07;
            16'd15004: data <= 8'hE0;
            16'd15005: data <= 8'h07;
            16'd15006: data <= 8'hE0;
            16'd15007: data <= 8'h07;
            16'd15008: data <= 8'hE0;
            16'd15009: data <= 8'h07;
            16'd15010: data <= 8'hE0;
            16'd15011: data <= 8'h07;
            16'd15012: data <= 8'hE0;
            16'd15013: data <= 8'h07;
            16'd15014: data <= 8'hE0;
            16'd15015: data <= 8'h07;
            16'd15016: data <= 8'hE0;
            16'd15017: data <= 8'h07;
            16'd15018: data <= 8'hE0;
            16'd15019: data <= 8'h07;
            16'd15020: data <= 8'hE0;
            16'd15021: data <= 8'h07;
            16'd15022: data <= 8'hE0;
            16'd15023: data <= 8'h07;
            16'd15024: data <= 8'hE0;
            16'd15025: data <= 8'h07;
            16'd15026: data <= 8'hE0;
            16'd15027: data <= 8'h07;
            16'd15028: data <= 8'hE0;
            16'd15029: data <= 8'h07;
            16'd15030: data <= 8'hE0;
            16'd15031: data <= 8'h07;
            16'd15032: data <= 8'hE0;
            16'd15033: data <= 8'h07;
            16'd15034: data <= 8'hE0;
            16'd15035: data <= 8'h07;
            16'd15036: data <= 8'hE0;
            16'd15037: data <= 8'h07;
            16'd15038: data <= 8'hE0;
            16'd15039: data <= 8'h07;
            16'd15040: data <= 8'hFF;
            16'd15041: data <= 8'hFF;
            16'd15042: data <= 8'hE0;
            16'd15043: data <= 8'h07;
            16'd15044: data <= 8'hE0;
            16'd15045: data <= 8'h07;
            16'd15046: data <= 8'hE0;
            16'd15047: data <= 8'h07;
            16'd15048: data <= 8'hE0;
            16'd15049: data <= 8'h07;
            16'd15050: data <= 8'hE0;
            16'd15051: data <= 8'h07;
            16'd15052: data <= 8'hE0;
            16'd15053: data <= 8'h07;
            16'd15054: data <= 8'hE0;
            16'd15055: data <= 8'h07;
            16'd15056: data <= 8'hE0;
            16'd15057: data <= 8'h07;
            16'd15058: data <= 8'hE0;
            16'd15059: data <= 8'h07;
            16'd15060: data <= 8'hE0;
            16'd15061: data <= 8'h07;
            16'd15062: data <= 8'hE0;
            16'd15063: data <= 8'h07;
            16'd15064: data <= 8'hE0;
            16'd15065: data <= 8'h07;
            16'd15066: data <= 8'hE0;
            16'd15067: data <= 8'h07;
            16'd15068: data <= 8'hE0;
            16'd15069: data <= 8'h07;
            16'd15070: data <= 8'hE0;
            16'd15071: data <= 8'h07;
            16'd15072: data <= 8'hE0;
            16'd15073: data <= 8'h07;
            16'd15074: data <= 8'hE0;
            16'd15075: data <= 8'h07;
            16'd15076: data <= 8'hE0;
            16'd15077: data <= 8'h07;
            16'd15078: data <= 8'hE0;
            16'd15079: data <= 8'h07;
            16'd15080: data <= 8'hFF;
            16'd15081: data <= 8'hFF;
            16'd15082: data <= 8'hE0;
            16'd15083: data <= 8'h07;
            16'd15084: data <= 8'hE0;
            16'd15085: data <= 8'h07;
            16'd15086: data <= 8'hE0;
            16'd15087: data <= 8'h07;
            16'd15088: data <= 8'hE0;
            16'd15089: data <= 8'h07;
            16'd15090: data <= 8'hE0;
            16'd15091: data <= 8'h07;
            16'd15092: data <= 8'hE0;
            16'd15093: data <= 8'h07;
            16'd15094: data <= 8'hE0;
            16'd15095: data <= 8'h07;
            16'd15096: data <= 8'hE0;
            16'd15097: data <= 8'h07;
            16'd15098: data <= 8'hE0;
            16'd15099: data <= 8'h07;
            16'd15100: data <= 8'hE0;
            16'd15101: data <= 8'h07;
            16'd15102: data <= 8'hE0;
            16'd15103: data <= 8'h07;
            16'd15104: data <= 8'hE0;
            16'd15105: data <= 8'h07;
            16'd15106: data <= 8'hE0;
            16'd15107: data <= 8'h07;
            16'd15108: data <= 8'hE0;
            16'd15109: data <= 8'h07;
            16'd15110: data <= 8'hE0;
            16'd15111: data <= 8'h07;
            16'd15112: data <= 8'hE0;
            16'd15113: data <= 8'h07;
            16'd15114: data <= 8'hE0;
            16'd15115: data <= 8'h07;
            16'd15116: data <= 8'hE0;
            16'd15117: data <= 8'h07;
            16'd15118: data <= 8'hE0;
            16'd15119: data <= 8'h07;
            16'd15120: data <= 8'hFF;
            16'd15121: data <= 8'hFF;
            16'd15122: data <= 8'hE0;
            16'd15123: data <= 8'h07;
            16'd15124: data <= 8'hE0;
            16'd15125: data <= 8'h07;
            16'd15126: data <= 8'hE0;
            16'd15127: data <= 8'h07;
            16'd15128: data <= 8'hE0;
            16'd15129: data <= 8'h07;
            16'd15130: data <= 8'hE0;
            16'd15131: data <= 8'h07;
            16'd15132: data <= 8'hE0;
            16'd15133: data <= 8'h07;
            16'd15134: data <= 8'hE0;
            16'd15135: data <= 8'h07;
            16'd15136: data <= 8'hE0;
            16'd15137: data <= 8'h07;
            16'd15138: data <= 8'hE0;
            16'd15139: data <= 8'h07;
            16'd15140: data <= 8'hE0;
            16'd15141: data <= 8'h07;
            16'd15142: data <= 8'hE0;
            16'd15143: data <= 8'h07;
            16'd15144: data <= 8'hE0;
            16'd15145: data <= 8'h07;
            16'd15146: data <= 8'hE0;
            16'd15147: data <= 8'h07;
            16'd15148: data <= 8'hE0;
            16'd15149: data <= 8'h07;
            16'd15150: data <= 8'hE0;
            16'd15151: data <= 8'h07;
            16'd15152: data <= 8'hE0;
            16'd15153: data <= 8'h07;
            16'd15154: data <= 8'hE0;
            16'd15155: data <= 8'h07;
            16'd15156: data <= 8'hE0;
            16'd15157: data <= 8'h07;
            16'd15158: data <= 8'hE0;
            16'd15159: data <= 8'h07;
            16'd15160: data <= 8'hFF;
            16'd15161: data <= 8'hFF;
            16'd15162: data <= 8'hE0;
            16'd15163: data <= 8'h07;
            16'd15164: data <= 8'hE0;
            16'd15165: data <= 8'h07;
            16'd15166: data <= 8'hE0;
            16'd15167: data <= 8'h07;
            16'd15168: data <= 8'hE0;
            16'd15169: data <= 8'h07;
            16'd15170: data <= 8'hE0;
            16'd15171: data <= 8'h07;
            16'd15172: data <= 8'hE0;
            16'd15173: data <= 8'h07;
            16'd15174: data <= 8'hE0;
            16'd15175: data <= 8'h07;
            16'd15176: data <= 8'hE0;
            16'd15177: data <= 8'h07;
            16'd15178: data <= 8'hE0;
            16'd15179: data <= 8'h07;
            16'd15180: data <= 8'hE0;
            16'd15181: data <= 8'h07;
            16'd15182: data <= 8'hE0;
            16'd15183: data <= 8'h07;
            16'd15184: data <= 8'hE0;
            16'd15185: data <= 8'h07;
            16'd15186: data <= 8'hE0;
            16'd15187: data <= 8'h07;
            16'd15188: data <= 8'hE0;
            16'd15189: data <= 8'h07;
            16'd15190: data <= 8'hE0;
            16'd15191: data <= 8'h07;
            16'd15192: data <= 8'hE0;
            16'd15193: data <= 8'h07;
            16'd15194: data <= 8'hE0;
            16'd15195: data <= 8'h07;
            16'd15196: data <= 8'hE0;
            16'd15197: data <= 8'h07;
            16'd15198: data <= 8'hE0;
            16'd15199: data <= 8'h07;
            16'd15200: data <= 8'hFF;
            16'd15201: data <= 8'hFF;
            16'd15202: data <= 8'hE0;
            16'd15203: data <= 8'h07;
            16'd15204: data <= 8'hE0;
            16'd15205: data <= 8'h07;
            16'd15206: data <= 8'hE0;
            16'd15207: data <= 8'h07;
            16'd15208: data <= 8'hE0;
            16'd15209: data <= 8'h07;
            16'd15210: data <= 8'hE0;
            16'd15211: data <= 8'h07;
            16'd15212: data <= 8'hE0;
            16'd15213: data <= 8'h07;
            16'd15214: data <= 8'hE0;
            16'd15215: data <= 8'h07;
            16'd15216: data <= 8'hE0;
            16'd15217: data <= 8'h07;
            16'd15218: data <= 8'hE0;
            16'd15219: data <= 8'h07;
            16'd15220: data <= 8'hE0;
            16'd15221: data <= 8'h07;
            16'd15222: data <= 8'hE0;
            16'd15223: data <= 8'h07;
            16'd15224: data <= 8'hE0;
            16'd15225: data <= 8'h07;
            16'd15226: data <= 8'hE0;
            16'd15227: data <= 8'h07;
            16'd15228: data <= 8'hE0;
            16'd15229: data <= 8'h07;
            16'd15230: data <= 8'hE0;
            16'd15231: data <= 8'h07;
            16'd15232: data <= 8'hE0;
            16'd15233: data <= 8'h07;
            16'd15234: data <= 8'hE0;
            16'd15235: data <= 8'h07;
            16'd15236: data <= 8'hE0;
            16'd15237: data <= 8'h07;
            16'd15238: data <= 8'hE0;
            16'd15239: data <= 8'h07;
            16'd15240: data <= 8'hFF;
            16'd15241: data <= 8'hFF;
            16'd15242: data <= 8'hE0;
            16'd15243: data <= 8'h07;
            16'd15244: data <= 8'hE0;
            16'd15245: data <= 8'h07;
            16'd15246: data <= 8'hE0;
            16'd15247: data <= 8'h07;
            16'd15248: data <= 8'hE0;
            16'd15249: data <= 8'h07;
            16'd15250: data <= 8'hE0;
            16'd15251: data <= 8'h07;
            16'd15252: data <= 8'hE0;
            16'd15253: data <= 8'h07;
            16'd15254: data <= 8'hE0;
            16'd15255: data <= 8'h07;
            16'd15256: data <= 8'hE0;
            16'd15257: data <= 8'h07;
            16'd15258: data <= 8'hE0;
            16'd15259: data <= 8'h07;
            16'd15260: data <= 8'hE0;
            16'd15261: data <= 8'h07;
            16'd15262: data <= 8'hE0;
            16'd15263: data <= 8'h07;
            16'd15264: data <= 8'hE0;
            16'd15265: data <= 8'h07;
            16'd15266: data <= 8'hE0;
            16'd15267: data <= 8'h07;
            16'd15268: data <= 8'hE0;
            16'd15269: data <= 8'h07;
            16'd15270: data <= 8'hE0;
            16'd15271: data <= 8'h07;
            16'd15272: data <= 8'hE0;
            16'd15273: data <= 8'h07;
            16'd15274: data <= 8'hE0;
            16'd15275: data <= 8'h07;
            16'd15276: data <= 8'hE0;
            16'd15277: data <= 8'h07;
            16'd15278: data <= 8'hE0;
            16'd15279: data <= 8'h07;
            16'd15280: data <= 8'hFF;
            16'd15281: data <= 8'hFF;
            16'd15282: data <= 8'hE0;
            16'd15283: data <= 8'h07;
            16'd15284: data <= 8'hE0;
            16'd15285: data <= 8'h07;
            16'd15286: data <= 8'hE0;
            16'd15287: data <= 8'h07;
            16'd15288: data <= 8'hE0;
            16'd15289: data <= 8'h07;
            16'd15290: data <= 8'hE0;
            16'd15291: data <= 8'h07;
            16'd15292: data <= 8'hE0;
            16'd15293: data <= 8'h07;
            16'd15294: data <= 8'hE0;
            16'd15295: data <= 8'h07;
            16'd15296: data <= 8'hE0;
            16'd15297: data <= 8'h07;
            16'd15298: data <= 8'hE0;
            16'd15299: data <= 8'h07;
            16'd15300: data <= 8'hE0;
            16'd15301: data <= 8'h07;
            16'd15302: data <= 8'hE0;
            16'd15303: data <= 8'h07;
            16'd15304: data <= 8'hE0;
            16'd15305: data <= 8'h07;
            16'd15306: data <= 8'hE0;
            16'd15307: data <= 8'h07;
            16'd15308: data <= 8'hE0;
            16'd15309: data <= 8'h07;
            16'd15310: data <= 8'hE0;
            16'd15311: data <= 8'h07;
            16'd15312: data <= 8'hE0;
            16'd15313: data <= 8'h07;
            16'd15314: data <= 8'hE0;
            16'd15315: data <= 8'h07;
            16'd15316: data <= 8'hE0;
            16'd15317: data <= 8'h07;
            16'd15318: data <= 8'hE0;
            16'd15319: data <= 8'h07;
            16'd15320: data <= 8'hFF;
            16'd15321: data <= 8'hFF;
            16'd15322: data <= 8'hE0;
            16'd15323: data <= 8'h07;
            16'd15324: data <= 8'hE0;
            16'd15325: data <= 8'h07;
            16'd15326: data <= 8'hE0;
            16'd15327: data <= 8'h07;
            16'd15328: data <= 8'hE0;
            16'd15329: data <= 8'h07;
            16'd15330: data <= 8'hE0;
            16'd15331: data <= 8'h07;
            16'd15332: data <= 8'hE0;
            16'd15333: data <= 8'h07;
            16'd15334: data <= 8'hE0;
            16'd15335: data <= 8'h07;
            16'd15336: data <= 8'hE0;
            16'd15337: data <= 8'h07;
            16'd15338: data <= 8'hE0;
            16'd15339: data <= 8'h07;
            16'd15340: data <= 8'hE0;
            16'd15341: data <= 8'h07;
            16'd15342: data <= 8'hE0;
            16'd15343: data <= 8'h07;
            16'd15344: data <= 8'hE0;
            16'd15345: data <= 8'h07;
            16'd15346: data <= 8'hE0;
            16'd15347: data <= 8'h07;
            16'd15348: data <= 8'hE0;
            16'd15349: data <= 8'h07;
            16'd15350: data <= 8'hE0;
            16'd15351: data <= 8'h07;
            16'd15352: data <= 8'hE0;
            16'd15353: data <= 8'h07;
            16'd15354: data <= 8'hE0;
            16'd15355: data <= 8'h07;
            16'd15356: data <= 8'hE0;
            16'd15357: data <= 8'h07;
            16'd15358: data <= 8'hE0;
            16'd15359: data <= 8'h07;
            16'd15360: data <= 8'hFF;
            16'd15361: data <= 8'hFF;
            16'd15362: data <= 8'hE0;
            16'd15363: data <= 8'h07;
            16'd15364: data <= 8'hE0;
            16'd15365: data <= 8'h07;
            16'd15366: data <= 8'hE0;
            16'd15367: data <= 8'h07;
            16'd15368: data <= 8'hE0;
            16'd15369: data <= 8'h07;
            16'd15370: data <= 8'hE0;
            16'd15371: data <= 8'h07;
            16'd15372: data <= 8'hE0;
            16'd15373: data <= 8'h07;
            16'd15374: data <= 8'hE0;
            16'd15375: data <= 8'h07;
            16'd15376: data <= 8'hE0;
            16'd15377: data <= 8'h07;
            16'd15378: data <= 8'hE0;
            16'd15379: data <= 8'h07;
            16'd15380: data <= 8'hE0;
            16'd15381: data <= 8'h07;
            16'd15382: data <= 8'hE0;
            16'd15383: data <= 8'h07;
            16'd15384: data <= 8'hE0;
            16'd15385: data <= 8'h07;
            16'd15386: data <= 8'hE0;
            16'd15387: data <= 8'h07;
            16'd15388: data <= 8'hE0;
            16'd15389: data <= 8'h07;
            16'd15390: data <= 8'hE0;
            16'd15391: data <= 8'h07;
            16'd15392: data <= 8'hE0;
            16'd15393: data <= 8'h07;
            16'd15394: data <= 8'hE0;
            16'd15395: data <= 8'h07;
            16'd15396: data <= 8'hE0;
            16'd15397: data <= 8'h07;
            16'd15398: data <= 8'hE0;
            16'd15399: data <= 8'h07;
            16'd15400: data <= 8'hFF;
            16'd15401: data <= 8'hFF;
            16'd15402: data <= 8'hE0;
            16'd15403: data <= 8'h07;
            16'd15404: data <= 8'hE0;
            16'd15405: data <= 8'h07;
            16'd15406: data <= 8'hE0;
            16'd15407: data <= 8'h07;
            16'd15408: data <= 8'hE0;
            16'd15409: data <= 8'h07;
            16'd15410: data <= 8'hE0;
            16'd15411: data <= 8'h07;
            16'd15412: data <= 8'hE0;
            16'd15413: data <= 8'h07;
            16'd15414: data <= 8'hE0;
            16'd15415: data <= 8'h07;
            16'd15416: data <= 8'hE0;
            16'd15417: data <= 8'h07;
            16'd15418: data <= 8'hE0;
            16'd15419: data <= 8'h07;
            16'd15420: data <= 8'hE0;
            16'd15421: data <= 8'h07;
            16'd15422: data <= 8'hE0;
            16'd15423: data <= 8'h07;
            16'd15424: data <= 8'hE0;
            16'd15425: data <= 8'h07;
            16'd15426: data <= 8'hE0;
            16'd15427: data <= 8'h07;
            16'd15428: data <= 8'hE0;
            16'd15429: data <= 8'h07;
            16'd15430: data <= 8'hE0;
            16'd15431: data <= 8'h07;
            16'd15432: data <= 8'hE0;
            16'd15433: data <= 8'h07;
            16'd15434: data <= 8'hE0;
            16'd15435: data <= 8'h07;
            16'd15436: data <= 8'hE0;
            16'd15437: data <= 8'h07;
            16'd15438: data <= 8'hE0;
            16'd15439: data <= 8'h07;
            16'd15440: data <= 8'hFF;
            16'd15441: data <= 8'hFF;
            16'd15442: data <= 8'hE0;
            16'd15443: data <= 8'h07;
            16'd15444: data <= 8'hE0;
            16'd15445: data <= 8'h07;
            16'd15446: data <= 8'hE0;
            16'd15447: data <= 8'h07;
            16'd15448: data <= 8'hE0;
            16'd15449: data <= 8'h07;
            16'd15450: data <= 8'hE0;
            16'd15451: data <= 8'h07;
            16'd15452: data <= 8'hE0;
            16'd15453: data <= 8'h07;
            16'd15454: data <= 8'hE0;
            16'd15455: data <= 8'h07;
            16'd15456: data <= 8'hE0;
            16'd15457: data <= 8'h07;
            16'd15458: data <= 8'hE0;
            16'd15459: data <= 8'h07;
            16'd15460: data <= 8'hE0;
            16'd15461: data <= 8'h07;
            16'd15462: data <= 8'hE0;
            16'd15463: data <= 8'h07;
            16'd15464: data <= 8'hE0;
            16'd15465: data <= 8'h07;
            16'd15466: data <= 8'hE0;
            16'd15467: data <= 8'h07;
            16'd15468: data <= 8'hE0;
            16'd15469: data <= 8'h07;
            16'd15470: data <= 8'hE0;
            16'd15471: data <= 8'h07;
            16'd15472: data <= 8'hE0;
            16'd15473: data <= 8'h07;
            16'd15474: data <= 8'hE0;
            16'd15475: data <= 8'h07;
            16'd15476: data <= 8'hE0;
            16'd15477: data <= 8'h07;
            16'd15478: data <= 8'hE0;
            16'd15479: data <= 8'h07;
            16'd15480: data <= 8'hFF;
            16'd15481: data <= 8'hFF;
            16'd15482: data <= 8'hE0;
            16'd15483: data <= 8'h07;
            16'd15484: data <= 8'hE0;
            16'd15485: data <= 8'h07;
            16'd15486: data <= 8'hE0;
            16'd15487: data <= 8'h07;
            16'd15488: data <= 8'hE0;
            16'd15489: data <= 8'h07;
            16'd15490: data <= 8'hE0;
            16'd15491: data <= 8'h07;
            16'd15492: data <= 8'hE0;
            16'd15493: data <= 8'h07;
            16'd15494: data <= 8'hE0;
            16'd15495: data <= 8'h07;
            16'd15496: data <= 8'hE0;
            16'd15497: data <= 8'h07;
            16'd15498: data <= 8'hE0;
            16'd15499: data <= 8'h07;
            16'd15500: data <= 8'hE0;
            16'd15501: data <= 8'h07;
            16'd15502: data <= 8'hE0;
            16'd15503: data <= 8'h07;
            16'd15504: data <= 8'hE0;
            16'd15505: data <= 8'h07;
            16'd15506: data <= 8'hE0;
            16'd15507: data <= 8'h07;
            16'd15508: data <= 8'hE0;
            16'd15509: data <= 8'h07;
            16'd15510: data <= 8'hE0;
            16'd15511: data <= 8'h07;
            16'd15512: data <= 8'hE0;
            16'd15513: data <= 8'h07;
            16'd15514: data <= 8'hE0;
            16'd15515: data <= 8'h07;
            16'd15516: data <= 8'hE0;
            16'd15517: data <= 8'h07;
            16'd15518: data <= 8'hE0;
            16'd15519: data <= 8'h07;
            16'd15520: data <= 8'hFF;
            16'd15521: data <= 8'hFF;
            16'd15522: data <= 8'hE0;
            16'd15523: data <= 8'h07;
            16'd15524: data <= 8'hE0;
            16'd15525: data <= 8'h07;
            16'd15526: data <= 8'hE0;
            16'd15527: data <= 8'h07;
            16'd15528: data <= 8'hE0;
            16'd15529: data <= 8'h07;
            16'd15530: data <= 8'hE0;
            16'd15531: data <= 8'h07;
            16'd15532: data <= 8'hE0;
            16'd15533: data <= 8'h07;
            16'd15534: data <= 8'hE0;
            16'd15535: data <= 8'h07;
            16'd15536: data <= 8'hE0;
            16'd15537: data <= 8'h07;
            16'd15538: data <= 8'hE0;
            16'd15539: data <= 8'h07;
            16'd15540: data <= 8'hE0;
            16'd15541: data <= 8'h07;
            16'd15542: data <= 8'hE0;
            16'd15543: data <= 8'h07;
            16'd15544: data <= 8'hE0;
            16'd15545: data <= 8'h07;
            16'd15546: data <= 8'hE0;
            16'd15547: data <= 8'h07;
            16'd15548: data <= 8'hE0;
            16'd15549: data <= 8'h07;
            16'd15550: data <= 8'hE0;
            16'd15551: data <= 8'h07;
            16'd15552: data <= 8'hE0;
            16'd15553: data <= 8'h07;
            16'd15554: data <= 8'hE0;
            16'd15555: data <= 8'h07;
            16'd15556: data <= 8'hE0;
            16'd15557: data <= 8'h07;
            16'd15558: data <= 8'hE0;
            16'd15559: data <= 8'h07;
            16'd15560: data <= 8'hFF;
            16'd15561: data <= 8'hFF;
            16'd15562: data <= 8'hE0;
            16'd15563: data <= 8'h07;
            16'd15564: data <= 8'hE0;
            16'd15565: data <= 8'h07;
            16'd15566: data <= 8'hE0;
            16'd15567: data <= 8'h07;
            16'd15568: data <= 8'hE0;
            16'd15569: data <= 8'h07;
            16'd15570: data <= 8'hE0;
            16'd15571: data <= 8'h07;
            16'd15572: data <= 8'hE0;
            16'd15573: data <= 8'h07;
            16'd15574: data <= 8'hE0;
            16'd15575: data <= 8'h07;
            16'd15576: data <= 8'hE0;
            16'd15577: data <= 8'h07;
            16'd15578: data <= 8'hE0;
            16'd15579: data <= 8'h07;
            16'd15580: data <= 8'hE0;
            16'd15581: data <= 8'h07;
            16'd15582: data <= 8'hE0;
            16'd15583: data <= 8'h07;
            16'd15584: data <= 8'hE0;
            16'd15585: data <= 8'h07;
            16'd15586: data <= 8'hE0;
            16'd15587: data <= 8'h07;
            16'd15588: data <= 8'hE0;
            16'd15589: data <= 8'h07;
            16'd15590: data <= 8'hE0;
            16'd15591: data <= 8'h07;
            16'd15592: data <= 8'hE0;
            16'd15593: data <= 8'h07;
            16'd15594: data <= 8'hE0;
            16'd15595: data <= 8'h07;
            16'd15596: data <= 8'hE0;
            16'd15597: data <= 8'h07;
            16'd15598: data <= 8'hE0;
            16'd15599: data <= 8'h07;
            16'd15600: data <= 8'hFF;
            16'd15601: data <= 8'hFF;
            16'd15602: data <= 8'hE0;
            16'd15603: data <= 8'h07;
            16'd15604: data <= 8'hE0;
            16'd15605: data <= 8'h07;
            16'd15606: data <= 8'hE0;
            16'd15607: data <= 8'h07;
            16'd15608: data <= 8'hE0;
            16'd15609: data <= 8'h07;
            16'd15610: data <= 8'hE0;
            16'd15611: data <= 8'h07;
            16'd15612: data <= 8'hE0;
            16'd15613: data <= 8'h07;
            16'd15614: data <= 8'hE0;
            16'd15615: data <= 8'h07;
            16'd15616: data <= 8'hE0;
            16'd15617: data <= 8'h07;
            16'd15618: data <= 8'hE0;
            16'd15619: data <= 8'h07;
            16'd15620: data <= 8'hE0;
            16'd15621: data <= 8'h07;
            16'd15622: data <= 8'hE0;
            16'd15623: data <= 8'h07;
            16'd15624: data <= 8'hE0;
            16'd15625: data <= 8'h07;
            16'd15626: data <= 8'hE0;
            16'd15627: data <= 8'h07;
            16'd15628: data <= 8'hE0;
            16'd15629: data <= 8'h07;
            16'd15630: data <= 8'hE0;
            16'd15631: data <= 8'h07;
            16'd15632: data <= 8'hE0;
            16'd15633: data <= 8'h07;
            16'd15634: data <= 8'hE0;
            16'd15635: data <= 8'h07;
            16'd15636: data <= 8'hE0;
            16'd15637: data <= 8'h07;
            16'd15638: data <= 8'hE0;
            16'd15639: data <= 8'h07;
            16'd15640: data <= 8'hFF;
            16'd15641: data <= 8'hFF;
            16'd15642: data <= 8'hE0;
            16'd15643: data <= 8'h07;
            16'd15644: data <= 8'hE0;
            16'd15645: data <= 8'h07;
            16'd15646: data <= 8'hE0;
            16'd15647: data <= 8'h07;
            16'd15648: data <= 8'hE0;
            16'd15649: data <= 8'h07;
            16'd15650: data <= 8'hE0;
            16'd15651: data <= 8'h07;
            16'd15652: data <= 8'hE0;
            16'd15653: data <= 8'h07;
            16'd15654: data <= 8'hE0;
            16'd15655: data <= 8'h07;
            16'd15656: data <= 8'hE0;
            16'd15657: data <= 8'h07;
            16'd15658: data <= 8'hE0;
            16'd15659: data <= 8'h07;
            16'd15660: data <= 8'hE0;
            16'd15661: data <= 8'h07;
            16'd15662: data <= 8'hE0;
            16'd15663: data <= 8'h07;
            16'd15664: data <= 8'hE0;
            16'd15665: data <= 8'h07;
            16'd15666: data <= 8'hE0;
            16'd15667: data <= 8'h07;
            16'd15668: data <= 8'hE0;
            16'd15669: data <= 8'h07;
            16'd15670: data <= 8'hE0;
            16'd15671: data <= 8'h07;
            16'd15672: data <= 8'hE0;
            16'd15673: data <= 8'h07;
            16'd15674: data <= 8'hE0;
            16'd15675: data <= 8'h07;
            16'd15676: data <= 8'hE0;
            16'd15677: data <= 8'h07;
            16'd15678: data <= 8'hE0;
            16'd15679: data <= 8'h07;
            16'd15680: data <= 8'hFF;
            16'd15681: data <= 8'hFF;
            16'd15682: data <= 8'hE0;
            16'd15683: data <= 8'h07;
            16'd15684: data <= 8'hE0;
            16'd15685: data <= 8'h07;
            16'd15686: data <= 8'hE0;
            16'd15687: data <= 8'h07;
            16'd15688: data <= 8'hE0;
            16'd15689: data <= 8'h07;
            16'd15690: data <= 8'hE0;
            16'd15691: data <= 8'h07;
            16'd15692: data <= 8'hE0;
            16'd15693: data <= 8'h07;
            16'd15694: data <= 8'hE0;
            16'd15695: data <= 8'h07;
            16'd15696: data <= 8'hE0;
            16'd15697: data <= 8'h07;
            16'd15698: data <= 8'hE0;
            16'd15699: data <= 8'h07;
            16'd15700: data <= 8'hE0;
            16'd15701: data <= 8'h07;
            16'd15702: data <= 8'hE0;
            16'd15703: data <= 8'h07;
            16'd15704: data <= 8'hE0;
            16'd15705: data <= 8'h07;
            16'd15706: data <= 8'hE0;
            16'd15707: data <= 8'h07;
            16'd15708: data <= 8'hE0;
            16'd15709: data <= 8'h07;
            16'd15710: data <= 8'hE0;
            16'd15711: data <= 8'h07;
            16'd15712: data <= 8'hE0;
            16'd15713: data <= 8'h07;
            16'd15714: data <= 8'hE0;
            16'd15715: data <= 8'h07;
            16'd15716: data <= 8'hE0;
            16'd15717: data <= 8'h07;
            16'd15718: data <= 8'hE0;
            16'd15719: data <= 8'h07;
            16'd15720: data <= 8'hFF;
            16'd15721: data <= 8'hFF;
            16'd15722: data <= 8'hE0;
            16'd15723: data <= 8'h07;
            16'd15724: data <= 8'hE0;
            16'd15725: data <= 8'h07;
            16'd15726: data <= 8'hE0;
            16'd15727: data <= 8'h07;
            16'd15728: data <= 8'hE0;
            16'd15729: data <= 8'h07;
            16'd15730: data <= 8'hE0;
            16'd15731: data <= 8'h07;
            16'd15732: data <= 8'hE0;
            16'd15733: data <= 8'h07;
            16'd15734: data <= 8'hE0;
            16'd15735: data <= 8'h07;
            16'd15736: data <= 8'hE0;
            16'd15737: data <= 8'h07;
            16'd15738: data <= 8'hE0;
            16'd15739: data <= 8'h07;
            16'd15740: data <= 8'hE0;
            16'd15741: data <= 8'h07;
            16'd15742: data <= 8'hE0;
            16'd15743: data <= 8'h07;
            16'd15744: data <= 8'hE0;
            16'd15745: data <= 8'h07;
            16'd15746: data <= 8'hE0;
            16'd15747: data <= 8'h07;
            16'd15748: data <= 8'hE0;
            16'd15749: data <= 8'h07;
            16'd15750: data <= 8'hE0;
            16'd15751: data <= 8'h07;
            16'd15752: data <= 8'hE0;
            16'd15753: data <= 8'h07;
            16'd15754: data <= 8'hE0;
            16'd15755: data <= 8'h07;
            16'd15756: data <= 8'hE0;
            16'd15757: data <= 8'h07;
            16'd15758: data <= 8'hE0;
            16'd15759: data <= 8'h07;
            16'd15760: data <= 8'hFF;
            16'd15761: data <= 8'hFF;
            16'd15762: data <= 8'hE0;
            16'd15763: data <= 8'h07;
            16'd15764: data <= 8'hE0;
            16'd15765: data <= 8'h07;
            16'd15766: data <= 8'hE0;
            16'd15767: data <= 8'h07;
            16'd15768: data <= 8'hE0;
            16'd15769: data <= 8'h07;
            16'd15770: data <= 8'hE0;
            16'd15771: data <= 8'h07;
            16'd15772: data <= 8'hE0;
            16'd15773: data <= 8'h07;
            16'd15774: data <= 8'hE0;
            16'd15775: data <= 8'h07;
            16'd15776: data <= 8'hE0;
            16'd15777: data <= 8'h07;
            16'd15778: data <= 8'hE0;
            16'd15779: data <= 8'h07;
            16'd15780: data <= 8'hE0;
            16'd15781: data <= 8'h07;
            16'd15782: data <= 8'hE0;
            16'd15783: data <= 8'h07;
            16'd15784: data <= 8'hE0;
            16'd15785: data <= 8'h07;
            16'd15786: data <= 8'hE0;
            16'd15787: data <= 8'h07;
            16'd15788: data <= 8'hE0;
            16'd15789: data <= 8'h07;
            16'd15790: data <= 8'hE0;
            16'd15791: data <= 8'h07;
            16'd15792: data <= 8'hE0;
            16'd15793: data <= 8'h07;
            16'd15794: data <= 8'hE0;
            16'd15795: data <= 8'h07;
            16'd15796: data <= 8'hE0;
            16'd15797: data <= 8'h07;
            16'd15798: data <= 8'hE0;
            16'd15799: data <= 8'h07;
            16'd15800: data <= 8'hFF;
            16'd15801: data <= 8'hFF;
            16'd15802: data <= 8'hE0;
            16'd15803: data <= 8'h07;
            16'd15804: data <= 8'hE0;
            16'd15805: data <= 8'h07;
            16'd15806: data <= 8'hE0;
            16'd15807: data <= 8'h07;
            16'd15808: data <= 8'hE0;
            16'd15809: data <= 8'h07;
            16'd15810: data <= 8'hE0;
            16'd15811: data <= 8'h07;
            16'd15812: data <= 8'hE0;
            16'd15813: data <= 8'h07;
            16'd15814: data <= 8'hE0;
            16'd15815: data <= 8'h07;
            16'd15816: data <= 8'hE0;
            16'd15817: data <= 8'h07;
            16'd15818: data <= 8'hE0;
            16'd15819: data <= 8'h07;
            16'd15820: data <= 8'hE0;
            16'd15821: data <= 8'h07;
            16'd15822: data <= 8'hE0;
            16'd15823: data <= 8'h07;
            16'd15824: data <= 8'hE0;
            16'd15825: data <= 8'h07;
            16'd15826: data <= 8'hE0;
            16'd15827: data <= 8'h07;
            16'd15828: data <= 8'hE0;
            16'd15829: data <= 8'h07;
            16'd15830: data <= 8'hE0;
            16'd15831: data <= 8'h07;
            16'd15832: data <= 8'hE0;
            16'd15833: data <= 8'h07;
            16'd15834: data <= 8'hE0;
            16'd15835: data <= 8'h07;
            16'd15836: data <= 8'hE0;
            16'd15837: data <= 8'h07;
            16'd15838: data <= 8'hE0;
            16'd15839: data <= 8'h07;
            16'd15840: data <= 8'hFF;
            16'd15841: data <= 8'hFF;
            16'd15842: data <= 8'hE0;
            16'd15843: data <= 8'h07;
            16'd15844: data <= 8'hE0;
            16'd15845: data <= 8'h07;
            16'd15846: data <= 8'hE0;
            16'd15847: data <= 8'h07;
            16'd15848: data <= 8'hE0;
            16'd15849: data <= 8'h07;
            16'd15850: data <= 8'hE0;
            16'd15851: data <= 8'h07;
            16'd15852: data <= 8'hE0;
            16'd15853: data <= 8'h07;
            16'd15854: data <= 8'hE0;
            16'd15855: data <= 8'h07;
            16'd15856: data <= 8'hE0;
            16'd15857: data <= 8'h07;
            16'd15858: data <= 8'hE0;
            16'd15859: data <= 8'h07;
            16'd15860: data <= 8'hE0;
            16'd15861: data <= 8'h07;
            16'd15862: data <= 8'hE0;
            16'd15863: data <= 8'h07;
            16'd15864: data <= 8'hE0;
            16'd15865: data <= 8'h07;
            16'd15866: data <= 8'hE0;
            16'd15867: data <= 8'h07;
            16'd15868: data <= 8'hE0;
            16'd15869: data <= 8'h07;
            16'd15870: data <= 8'hE0;
            16'd15871: data <= 8'h07;
            16'd15872: data <= 8'hE0;
            16'd15873: data <= 8'h07;
            16'd15874: data <= 8'hE0;
            16'd15875: data <= 8'h07;
            16'd15876: data <= 8'hE0;
            16'd15877: data <= 8'h07;
            16'd15878: data <= 8'hE0;
            16'd15879: data <= 8'h07;
            16'd15880: data <= 8'hFF;
            16'd15881: data <= 8'hFF;
            16'd15882: data <= 8'hE0;
            16'd15883: data <= 8'h07;
            16'd15884: data <= 8'hE0;
            16'd15885: data <= 8'h07;
            16'd15886: data <= 8'hE0;
            16'd15887: data <= 8'h07;
            16'd15888: data <= 8'hE0;
            16'd15889: data <= 8'h07;
            16'd15890: data <= 8'hE0;
            16'd15891: data <= 8'h07;
            16'd15892: data <= 8'hE0;
            16'd15893: data <= 8'h07;
            16'd15894: data <= 8'hE0;
            16'd15895: data <= 8'h07;
            16'd15896: data <= 8'hE0;
            16'd15897: data <= 8'h07;
            16'd15898: data <= 8'hE0;
            16'd15899: data <= 8'h07;
            16'd15900: data <= 8'hE0;
            16'd15901: data <= 8'h07;
            16'd15902: data <= 8'hE0;
            16'd15903: data <= 8'h07;
            16'd15904: data <= 8'hE0;
            16'd15905: data <= 8'h07;
            16'd15906: data <= 8'hE0;
            16'd15907: data <= 8'h07;
            16'd15908: data <= 8'hE0;
            16'd15909: data <= 8'h07;
            16'd15910: data <= 8'hE0;
            16'd15911: data <= 8'h07;
            16'd15912: data <= 8'hE0;
            16'd15913: data <= 8'h07;
            16'd15914: data <= 8'hE0;
            16'd15915: data <= 8'h07;
            16'd15916: data <= 8'hE0;
            16'd15917: data <= 8'h07;
            16'd15918: data <= 8'hE0;
            16'd15919: data <= 8'h07;
            16'd15920: data <= 8'hFF;
            16'd15921: data <= 8'hFF;
            16'd15922: data <= 8'hE0;
            16'd15923: data <= 8'h07;
            16'd15924: data <= 8'hE0;
            16'd15925: data <= 8'h07;
            16'd15926: data <= 8'hE0;
            16'd15927: data <= 8'h07;
            16'd15928: data <= 8'hE0;
            16'd15929: data <= 8'h07;
            16'd15930: data <= 8'hE0;
            16'd15931: data <= 8'h07;
            16'd15932: data <= 8'hE0;
            16'd15933: data <= 8'h07;
            16'd15934: data <= 8'hE0;
            16'd15935: data <= 8'h07;
            16'd15936: data <= 8'hE0;
            16'd15937: data <= 8'h07;
            16'd15938: data <= 8'hE0;
            16'd15939: data <= 8'h07;
            16'd15940: data <= 8'hE0;
            16'd15941: data <= 8'h07;
            16'd15942: data <= 8'hE0;
            16'd15943: data <= 8'h07;
            16'd15944: data <= 8'hE0;
            16'd15945: data <= 8'h07;
            16'd15946: data <= 8'hE0;
            16'd15947: data <= 8'h07;
            16'd15948: data <= 8'hE0;
            16'd15949: data <= 8'h07;
            16'd15950: data <= 8'hE0;
            16'd15951: data <= 8'h07;
            16'd15952: data <= 8'hE0;
            16'd15953: data <= 8'h07;
            16'd15954: data <= 8'hE0;
            16'd15955: data <= 8'h07;
            16'd15956: data <= 8'hE0;
            16'd15957: data <= 8'h07;
            16'd15958: data <= 8'hE0;
            16'd15959: data <= 8'h07;
            16'd15960: data <= 8'hFF;
            16'd15961: data <= 8'hFF;
            16'd15962: data <= 8'hE0;
            16'd15963: data <= 8'h07;
            16'd15964: data <= 8'hE0;
            16'd15965: data <= 8'h07;
            16'd15966: data <= 8'hE0;
            16'd15967: data <= 8'h07;
            16'd15968: data <= 8'hE0;
            16'd15969: data <= 8'h07;
            16'd15970: data <= 8'hE0;
            16'd15971: data <= 8'h07;
            16'd15972: data <= 8'hE0;
            16'd15973: data <= 8'h07;
            16'd15974: data <= 8'hE0;
            16'd15975: data <= 8'h07;
            16'd15976: data <= 8'hE0;
            16'd15977: data <= 8'h07;
            16'd15978: data <= 8'hE0;
            16'd15979: data <= 8'h07;
            16'd15980: data <= 8'hE0;
            16'd15981: data <= 8'h07;
            16'd15982: data <= 8'hE0;
            16'd15983: data <= 8'h07;
            16'd15984: data <= 8'hE0;
            16'd15985: data <= 8'h07;
            16'd15986: data <= 8'hE0;
            16'd15987: data <= 8'h07;
            16'd15988: data <= 8'hE0;
            16'd15989: data <= 8'h07;
            16'd15990: data <= 8'hE0;
            16'd15991: data <= 8'h07;
            16'd15992: data <= 8'hE0;
            16'd15993: data <= 8'h07;
            16'd15994: data <= 8'hE0;
            16'd15995: data <= 8'h07;
            16'd15996: data <= 8'hE0;
            16'd15997: data <= 8'h07;
            16'd15998: data <= 8'hE0;
            16'd15999: data <= 8'h07;
            16'd16000: data <= 8'hFF;
            16'd16001: data <= 8'hFF;
            16'd16002: data <= 8'hE0;
            16'd16003: data <= 8'h07;
            16'd16004: data <= 8'hE0;
            16'd16005: data <= 8'h07;
            16'd16006: data <= 8'hE0;
            16'd16007: data <= 8'h07;
            16'd16008: data <= 8'hE0;
            16'd16009: data <= 8'h07;
            16'd16010: data <= 8'hE0;
            16'd16011: data <= 8'h07;
            16'd16012: data <= 8'hE0;
            16'd16013: data <= 8'h07;
            16'd16014: data <= 8'hE0;
            16'd16015: data <= 8'h07;
            16'd16016: data <= 8'hE0;
            16'd16017: data <= 8'h07;
            16'd16018: data <= 8'hE0;
            16'd16019: data <= 8'h07;
            16'd16020: data <= 8'hE0;
            16'd16021: data <= 8'h07;
            16'd16022: data <= 8'hE0;
            16'd16023: data <= 8'h07;
            16'd16024: data <= 8'hE0;
            16'd16025: data <= 8'h07;
            16'd16026: data <= 8'hE0;
            16'd16027: data <= 8'h07;
            16'd16028: data <= 8'hE0;
            16'd16029: data <= 8'h07;
            16'd16030: data <= 8'hE0;
            16'd16031: data <= 8'h07;
            16'd16032: data <= 8'hE0;
            16'd16033: data <= 8'h07;
            16'd16034: data <= 8'hE0;
            16'd16035: data <= 8'h07;
            16'd16036: data <= 8'hE0;
            16'd16037: data <= 8'h07;
            16'd16038: data <= 8'hE0;
            16'd16039: data <= 8'h07;
            16'd16040: data <= 8'hFF;
            16'd16041: data <= 8'hFF;
            16'd16042: data <= 8'hE0;
            16'd16043: data <= 8'h07;
            16'd16044: data <= 8'hE0;
            16'd16045: data <= 8'h07;
            16'd16046: data <= 8'hE0;
            16'd16047: data <= 8'h07;
            16'd16048: data <= 8'hE0;
            16'd16049: data <= 8'h07;
            16'd16050: data <= 8'hE0;
            16'd16051: data <= 8'h07;
            16'd16052: data <= 8'hE0;
            16'd16053: data <= 8'h07;
            16'd16054: data <= 8'hE0;
            16'd16055: data <= 8'h07;
            16'd16056: data <= 8'hE0;
            16'd16057: data <= 8'h07;
            16'd16058: data <= 8'hE0;
            16'd16059: data <= 8'h07;
            16'd16060: data <= 8'hE0;
            16'd16061: data <= 8'h07;
            16'd16062: data <= 8'hE0;
            16'd16063: data <= 8'h07;
            16'd16064: data <= 8'hE0;
            16'd16065: data <= 8'h07;
            16'd16066: data <= 8'hE0;
            16'd16067: data <= 8'h07;
            16'd16068: data <= 8'hE0;
            16'd16069: data <= 8'h07;
            16'd16070: data <= 8'hE0;
            16'd16071: data <= 8'h07;
            16'd16072: data <= 8'hE0;
            16'd16073: data <= 8'h07;
            16'd16074: data <= 8'hE0;
            16'd16075: data <= 8'h07;
            16'd16076: data <= 8'hE0;
            16'd16077: data <= 8'h07;
            16'd16078: data <= 8'hE0;
            16'd16079: data <= 8'h07;
            16'd16080: data <= 8'hFF;
            16'd16081: data <= 8'hFF;
            16'd16082: data <= 8'hE0;
            16'd16083: data <= 8'h07;
            16'd16084: data <= 8'hE0;
            16'd16085: data <= 8'h07;
            16'd16086: data <= 8'hE0;
            16'd16087: data <= 8'h07;
            16'd16088: data <= 8'hE0;
            16'd16089: data <= 8'h07;
            16'd16090: data <= 8'hE0;
            16'd16091: data <= 8'h07;
            16'd16092: data <= 8'hE0;
            16'd16093: data <= 8'h07;
            16'd16094: data <= 8'hE0;
            16'd16095: data <= 8'h07;
            16'd16096: data <= 8'hE0;
            16'd16097: data <= 8'h07;
            16'd16098: data <= 8'hE0;
            16'd16099: data <= 8'h07;
            16'd16100: data <= 8'hE0;
            16'd16101: data <= 8'h07;
            16'd16102: data <= 8'hE0;
            16'd16103: data <= 8'h07;
            16'd16104: data <= 8'hE0;
            16'd16105: data <= 8'h07;
            16'd16106: data <= 8'hE0;
            16'd16107: data <= 8'h07;
            16'd16108: data <= 8'hE0;
            16'd16109: data <= 8'h07;
            16'd16110: data <= 8'hE0;
            16'd16111: data <= 8'h07;
            16'd16112: data <= 8'hE0;
            16'd16113: data <= 8'h07;
            16'd16114: data <= 8'hE0;
            16'd16115: data <= 8'h07;
            16'd16116: data <= 8'hE0;
            16'd16117: data <= 8'h07;
            16'd16118: data <= 8'hE0;
            16'd16119: data <= 8'h07;
            16'd16120: data <= 8'hFF;
            16'd16121: data <= 8'hFF;
            16'd16122: data <= 8'hE0;
            16'd16123: data <= 8'h07;
            16'd16124: data <= 8'hE0;
            16'd16125: data <= 8'h07;
            16'd16126: data <= 8'hE0;
            16'd16127: data <= 8'h07;
            16'd16128: data <= 8'hE0;
            16'd16129: data <= 8'h07;
            16'd16130: data <= 8'hE0;
            16'd16131: data <= 8'h07;
            16'd16132: data <= 8'hE0;
            16'd16133: data <= 8'h07;
            16'd16134: data <= 8'hE0;
            16'd16135: data <= 8'h07;
            16'd16136: data <= 8'hE0;
            16'd16137: data <= 8'h07;
            16'd16138: data <= 8'hE0;
            16'd16139: data <= 8'h07;
            16'd16140: data <= 8'hE0;
            16'd16141: data <= 8'h07;
            16'd16142: data <= 8'hE0;
            16'd16143: data <= 8'h07;
            16'd16144: data <= 8'hE0;
            16'd16145: data <= 8'h07;
            16'd16146: data <= 8'hE0;
            16'd16147: data <= 8'h07;
            16'd16148: data <= 8'hE0;
            16'd16149: data <= 8'h07;
            16'd16150: data <= 8'hE0;
            16'd16151: data <= 8'h07;
            16'd16152: data <= 8'hE0;
            16'd16153: data <= 8'h07;
            16'd16154: data <= 8'hE0;
            16'd16155: data <= 8'h07;
            16'd16156: data <= 8'hE0;
            16'd16157: data <= 8'h07;
            16'd16158: data <= 8'hE0;
            16'd16159: data <= 8'h07;
            16'd16160: data <= 8'hFF;
            16'd16161: data <= 8'hFF;
            16'd16162: data <= 8'hE0;
            16'd16163: data <= 8'h07;
            16'd16164: data <= 8'hE0;
            16'd16165: data <= 8'h07;
            16'd16166: data <= 8'hE0;
            16'd16167: data <= 8'h07;
            16'd16168: data <= 8'hE0;
            16'd16169: data <= 8'h07;
            16'd16170: data <= 8'hE0;
            16'd16171: data <= 8'h07;
            16'd16172: data <= 8'hE0;
            16'd16173: data <= 8'h07;
            16'd16174: data <= 8'hE0;
            16'd16175: data <= 8'h07;
            16'd16176: data <= 8'hE0;
            16'd16177: data <= 8'h07;
            16'd16178: data <= 8'hE0;
            16'd16179: data <= 8'h07;
            16'd16180: data <= 8'hE0;
            16'd16181: data <= 8'h07;
            16'd16182: data <= 8'hE0;
            16'd16183: data <= 8'h07;
            16'd16184: data <= 8'hE0;
            16'd16185: data <= 8'h07;
            16'd16186: data <= 8'hE0;
            16'd16187: data <= 8'h07;
            16'd16188: data <= 8'hE0;
            16'd16189: data <= 8'h07;
            16'd16190: data <= 8'hE0;
            16'd16191: data <= 8'h07;
            16'd16192: data <= 8'hE0;
            16'd16193: data <= 8'h07;
            16'd16194: data <= 8'hE0;
            16'd16195: data <= 8'h07;
            16'd16196: data <= 8'hE0;
            16'd16197: data <= 8'h07;
            16'd16198: data <= 8'hE0;
            16'd16199: data <= 8'h07;
            16'd16200: data <= 8'hFF;
            16'd16201: data <= 8'hFF;
            16'd16202: data <= 8'hE0;
            16'd16203: data <= 8'h07;
            16'd16204: data <= 8'hE0;
            16'd16205: data <= 8'h07;
            16'd16206: data <= 8'hE0;
            16'd16207: data <= 8'h07;
            16'd16208: data <= 8'hE0;
            16'd16209: data <= 8'h07;
            16'd16210: data <= 8'hE0;
            16'd16211: data <= 8'h07;
            16'd16212: data <= 8'hE0;
            16'd16213: data <= 8'h07;
            16'd16214: data <= 8'hE0;
            16'd16215: data <= 8'h07;
            16'd16216: data <= 8'hE0;
            16'd16217: data <= 8'h07;
            16'd16218: data <= 8'hE0;
            16'd16219: data <= 8'h07;
            16'd16220: data <= 8'hE0;
            16'd16221: data <= 8'h07;
            16'd16222: data <= 8'hE0;
            16'd16223: data <= 8'h07;
            16'd16224: data <= 8'hE0;
            16'd16225: data <= 8'h07;
            16'd16226: data <= 8'hE0;
            16'd16227: data <= 8'h07;
            16'd16228: data <= 8'hE0;
            16'd16229: data <= 8'h07;
            16'd16230: data <= 8'hE0;
            16'd16231: data <= 8'h07;
            16'd16232: data <= 8'hE0;
            16'd16233: data <= 8'h07;
            16'd16234: data <= 8'hE0;
            16'd16235: data <= 8'h07;
            16'd16236: data <= 8'hE0;
            16'd16237: data <= 8'h07;
            16'd16238: data <= 8'hE0;
            16'd16239: data <= 8'h07;
            16'd16240: data <= 8'hFF;
            16'd16241: data <= 8'hFF;
            16'd16242: data <= 8'hE0;
            16'd16243: data <= 8'h07;
            16'd16244: data <= 8'hE0;
            16'd16245: data <= 8'h07;
            16'd16246: data <= 8'hE0;
            16'd16247: data <= 8'h07;
            16'd16248: data <= 8'hE0;
            16'd16249: data <= 8'h07;
            16'd16250: data <= 8'hE0;
            16'd16251: data <= 8'h07;
            16'd16252: data <= 8'hE0;
            16'd16253: data <= 8'h07;
            16'd16254: data <= 8'hE0;
            16'd16255: data <= 8'h07;
            16'd16256: data <= 8'hE0;
            16'd16257: data <= 8'h07;
            16'd16258: data <= 8'hE0;
            16'd16259: data <= 8'h07;
            16'd16260: data <= 8'hE0;
            16'd16261: data <= 8'h07;
            16'd16262: data <= 8'hE0;
            16'd16263: data <= 8'h07;
            16'd16264: data <= 8'hE0;
            16'd16265: data <= 8'h07;
            16'd16266: data <= 8'hE0;
            16'd16267: data <= 8'h07;
            16'd16268: data <= 8'hE0;
            16'd16269: data <= 8'h07;
            16'd16270: data <= 8'hE0;
            16'd16271: data <= 8'h07;
            16'd16272: data <= 8'hE0;
            16'd16273: data <= 8'h07;
            16'd16274: data <= 8'hE0;
            16'd16275: data <= 8'h07;
            16'd16276: data <= 8'hE0;
            16'd16277: data <= 8'h07;
            16'd16278: data <= 8'hE0;
            16'd16279: data <= 8'h07;
            16'd16280: data <= 8'hFF;
            16'd16281: data <= 8'hFF;
            16'd16282: data <= 8'hE0;
            16'd16283: data <= 8'h07;
            16'd16284: data <= 8'hE0;
            16'd16285: data <= 8'h07;
            16'd16286: data <= 8'hE0;
            16'd16287: data <= 8'h07;
            16'd16288: data <= 8'hE0;
            16'd16289: data <= 8'h07;
            16'd16290: data <= 8'hE0;
            16'd16291: data <= 8'h07;
            16'd16292: data <= 8'hE0;
            16'd16293: data <= 8'h07;
            16'd16294: data <= 8'hE0;
            16'd16295: data <= 8'h07;
            16'd16296: data <= 8'hE0;
            16'd16297: data <= 8'h07;
            16'd16298: data <= 8'hE0;
            16'd16299: data <= 8'h07;
            16'd16300: data <= 8'hE0;
            16'd16301: data <= 8'h07;
            16'd16302: data <= 8'hE0;
            16'd16303: data <= 8'h07;
            16'd16304: data <= 8'hE0;
            16'd16305: data <= 8'h07;
            16'd16306: data <= 8'hE0;
            16'd16307: data <= 8'h07;
            16'd16308: data <= 8'hE0;
            16'd16309: data <= 8'h07;
            16'd16310: data <= 8'hE0;
            16'd16311: data <= 8'h07;
            16'd16312: data <= 8'hE0;
            16'd16313: data <= 8'h07;
            16'd16314: data <= 8'hE0;
            16'd16315: data <= 8'h07;
            16'd16316: data <= 8'hE0;
            16'd16317: data <= 8'h07;
            16'd16318: data <= 8'hE0;
            16'd16319: data <= 8'h07;
            16'd16320: data <= 8'hFF;
            16'd16321: data <= 8'hFF;
            16'd16322: data <= 8'hE0;
            16'd16323: data <= 8'h07;
            16'd16324: data <= 8'hE0;
            16'd16325: data <= 8'h07;
            16'd16326: data <= 8'hE0;
            16'd16327: data <= 8'h07;
            16'd16328: data <= 8'hE0;
            16'd16329: data <= 8'h07;
            16'd16330: data <= 8'hE0;
            16'd16331: data <= 8'h07;
            16'd16332: data <= 8'hE0;
            16'd16333: data <= 8'h07;
            16'd16334: data <= 8'hE0;
            16'd16335: data <= 8'h07;
            16'd16336: data <= 8'hE0;
            16'd16337: data <= 8'h07;
            16'd16338: data <= 8'hE0;
            16'd16339: data <= 8'h07;
            16'd16340: data <= 8'hE0;
            16'd16341: data <= 8'h07;
            16'd16342: data <= 8'hE0;
            16'd16343: data <= 8'h07;
            16'd16344: data <= 8'hE0;
            16'd16345: data <= 8'h07;
            16'd16346: data <= 8'hE0;
            16'd16347: data <= 8'h07;
            16'd16348: data <= 8'hE0;
            16'd16349: data <= 8'h07;
            16'd16350: data <= 8'hE0;
            16'd16351: data <= 8'h07;
            16'd16352: data <= 8'hE0;
            16'd16353: data <= 8'h07;
            16'd16354: data <= 8'hE0;
            16'd16355: data <= 8'h07;
            16'd16356: data <= 8'hE0;
            16'd16357: data <= 8'h07;
            16'd16358: data <= 8'hE0;
            16'd16359: data <= 8'h07;
            16'd16360: data <= 8'hFF;
            16'd16361: data <= 8'hFF;
            16'd16362: data <= 8'hE0;
            16'd16363: data <= 8'h07;
            16'd16364: data <= 8'hE0;
            16'd16365: data <= 8'h07;
            16'd16366: data <= 8'hE0;
            16'd16367: data <= 8'h07;
            16'd16368: data <= 8'hE0;
            16'd16369: data <= 8'h07;
            16'd16370: data <= 8'hE0;
            16'd16371: data <= 8'h07;
            16'd16372: data <= 8'hE0;
            16'd16373: data <= 8'h07;
            16'd16374: data <= 8'hE0;
            16'd16375: data <= 8'h07;
            16'd16376: data <= 8'hE0;
            16'd16377: data <= 8'h07;
            16'd16378: data <= 8'hE0;
            16'd16379: data <= 8'h07;
            16'd16380: data <= 8'hE0;
            16'd16381: data <= 8'h07;
            16'd16382: data <= 8'hE0;
            16'd16383: data <= 8'h07;
            16'd16384: data <= 8'hE0;
            16'd16385: data <= 8'h07;
            16'd16386: data <= 8'hE0;
            16'd16387: data <= 8'h07;
            16'd16388: data <= 8'hE0;
            16'd16389: data <= 8'h07;
            16'd16390: data <= 8'hE0;
            16'd16391: data <= 8'h07;
            16'd16392: data <= 8'hE0;
            16'd16393: data <= 8'h07;
            16'd16394: data <= 8'hE0;
            16'd16395: data <= 8'h07;
            16'd16396: data <= 8'hE0;
            16'd16397: data <= 8'h07;
            16'd16398: data <= 8'hE0;
            16'd16399: data <= 8'h07;
            16'd16400: data <= 8'hFF;
            16'd16401: data <= 8'hFF;
            16'd16402: data <= 8'hE0;
            16'd16403: data <= 8'h07;
            16'd16404: data <= 8'hE0;
            16'd16405: data <= 8'h07;
            16'd16406: data <= 8'hE0;
            16'd16407: data <= 8'h07;
            16'd16408: data <= 8'hE0;
            16'd16409: data <= 8'h07;
            16'd16410: data <= 8'hE0;
            16'd16411: data <= 8'h07;
            16'd16412: data <= 8'hE0;
            16'd16413: data <= 8'h07;
            16'd16414: data <= 8'hE0;
            16'd16415: data <= 8'h07;
            16'd16416: data <= 8'hE0;
            16'd16417: data <= 8'h07;
            16'd16418: data <= 8'hE0;
            16'd16419: data <= 8'h07;
            16'd16420: data <= 8'hE0;
            16'd16421: data <= 8'h07;
            16'd16422: data <= 8'hE0;
            16'd16423: data <= 8'h07;
            16'd16424: data <= 8'hE0;
            16'd16425: data <= 8'h07;
            16'd16426: data <= 8'hE0;
            16'd16427: data <= 8'h07;
            16'd16428: data <= 8'hE0;
            16'd16429: data <= 8'h07;
            16'd16430: data <= 8'hE0;
            16'd16431: data <= 8'h07;
            16'd16432: data <= 8'hE0;
            16'd16433: data <= 8'h07;
            16'd16434: data <= 8'hE0;
            16'd16435: data <= 8'h07;
            16'd16436: data <= 8'hE0;
            16'd16437: data <= 8'h07;
            16'd16438: data <= 8'hE0;
            16'd16439: data <= 8'h07;
            16'd16440: data <= 8'hFF;
            16'd16441: data <= 8'hFF;
            16'd16442: data <= 8'hE0;
            16'd16443: data <= 8'h07;
            16'd16444: data <= 8'hE0;
            16'd16445: data <= 8'h07;
            16'd16446: data <= 8'hE0;
            16'd16447: data <= 8'h07;
            16'd16448: data <= 8'hE0;
            16'd16449: data <= 8'h07;
            16'd16450: data <= 8'hE0;
            16'd16451: data <= 8'h07;
            16'd16452: data <= 8'hE0;
            16'd16453: data <= 8'h07;
            16'd16454: data <= 8'hE0;
            16'd16455: data <= 8'h07;
            16'd16456: data <= 8'hE0;
            16'd16457: data <= 8'h07;
            16'd16458: data <= 8'hE0;
            16'd16459: data <= 8'h07;
            16'd16460: data <= 8'hE0;
            16'd16461: data <= 8'h07;
            16'd16462: data <= 8'hE0;
            16'd16463: data <= 8'h07;
            16'd16464: data <= 8'hE0;
            16'd16465: data <= 8'h07;
            16'd16466: data <= 8'hE0;
            16'd16467: data <= 8'h07;
            16'd16468: data <= 8'hE0;
            16'd16469: data <= 8'h07;
            16'd16470: data <= 8'hE0;
            16'd16471: data <= 8'h07;
            16'd16472: data <= 8'hE0;
            16'd16473: data <= 8'h07;
            16'd16474: data <= 8'hE0;
            16'd16475: data <= 8'h07;
            16'd16476: data <= 8'hE0;
            16'd16477: data <= 8'h07;
            16'd16478: data <= 8'hE0;
            16'd16479: data <= 8'h07;
            16'd16480: data <= 8'hFF;
            16'd16481: data <= 8'hFF;
            16'd16482: data <= 8'hE0;
            16'd16483: data <= 8'h07;
            16'd16484: data <= 8'hE0;
            16'd16485: data <= 8'h07;
            16'd16486: data <= 8'hE0;
            16'd16487: data <= 8'h07;
            16'd16488: data <= 8'hE0;
            16'd16489: data <= 8'h07;
            16'd16490: data <= 8'hE0;
            16'd16491: data <= 8'h07;
            16'd16492: data <= 8'hE0;
            16'd16493: data <= 8'h07;
            16'd16494: data <= 8'hE0;
            16'd16495: data <= 8'h07;
            16'd16496: data <= 8'hE0;
            16'd16497: data <= 8'h07;
            16'd16498: data <= 8'hE0;
            16'd16499: data <= 8'h07;
            16'd16500: data <= 8'hE0;
            16'd16501: data <= 8'h07;
            16'd16502: data <= 8'hE0;
            16'd16503: data <= 8'h07;
            16'd16504: data <= 8'hE0;
            16'd16505: data <= 8'h07;
            16'd16506: data <= 8'hE0;
            16'd16507: data <= 8'h07;
            16'd16508: data <= 8'hE0;
            16'd16509: data <= 8'h07;
            16'd16510: data <= 8'hE0;
            16'd16511: data <= 8'h07;
            16'd16512: data <= 8'hE0;
            16'd16513: data <= 8'h07;
            16'd16514: data <= 8'hE0;
            16'd16515: data <= 8'h07;
            16'd16516: data <= 8'hE0;
            16'd16517: data <= 8'h07;
            16'd16518: data <= 8'hE0;
            16'd16519: data <= 8'h07;
            16'd16520: data <= 8'hFF;
            16'd16521: data <= 8'hFF;
            16'd16522: data <= 8'hE0;
            16'd16523: data <= 8'h07;
            16'd16524: data <= 8'hE0;
            16'd16525: data <= 8'h07;
            16'd16526: data <= 8'hE0;
            16'd16527: data <= 8'h07;
            16'd16528: data <= 8'hE0;
            16'd16529: data <= 8'h07;
            16'd16530: data <= 8'hE0;
            16'd16531: data <= 8'h07;
            16'd16532: data <= 8'hE0;
            16'd16533: data <= 8'h07;
            16'd16534: data <= 8'hE0;
            16'd16535: data <= 8'h07;
            16'd16536: data <= 8'hE0;
            16'd16537: data <= 8'h07;
            16'd16538: data <= 8'hE0;
            16'd16539: data <= 8'h07;
            16'd16540: data <= 8'hE0;
            16'd16541: data <= 8'h07;
            16'd16542: data <= 8'hE0;
            16'd16543: data <= 8'h07;
            16'd16544: data <= 8'hE0;
            16'd16545: data <= 8'h07;
            16'd16546: data <= 8'hE0;
            16'd16547: data <= 8'h07;
            16'd16548: data <= 8'hE0;
            16'd16549: data <= 8'h07;
            16'd16550: data <= 8'hE0;
            16'd16551: data <= 8'h07;
            16'd16552: data <= 8'hE0;
            16'd16553: data <= 8'h07;
            16'd16554: data <= 8'hE0;
            16'd16555: data <= 8'h07;
            16'd16556: data <= 8'hE0;
            16'd16557: data <= 8'h07;
            16'd16558: data <= 8'hE0;
            16'd16559: data <= 8'h07;
            16'd16560: data <= 8'hFF;
            16'd16561: data <= 8'hFF;
            16'd16562: data <= 8'hE0;
            16'd16563: data <= 8'h07;
            16'd16564: data <= 8'hE0;
            16'd16565: data <= 8'h07;
            16'd16566: data <= 8'hE0;
            16'd16567: data <= 8'h07;
            16'd16568: data <= 8'hE0;
            16'd16569: data <= 8'h07;
            16'd16570: data <= 8'hE0;
            16'd16571: data <= 8'h07;
            16'd16572: data <= 8'hE0;
            16'd16573: data <= 8'h07;
            16'd16574: data <= 8'hE0;
            16'd16575: data <= 8'h07;
            16'd16576: data <= 8'hE0;
            16'd16577: data <= 8'h07;
            16'd16578: data <= 8'hE0;
            16'd16579: data <= 8'h07;
            16'd16580: data <= 8'hE0;
            16'd16581: data <= 8'h07;
            16'd16582: data <= 8'hE0;
            16'd16583: data <= 8'h07;
            16'd16584: data <= 8'hE0;
            16'd16585: data <= 8'h07;
            16'd16586: data <= 8'hE0;
            16'd16587: data <= 8'h07;
            16'd16588: data <= 8'hE0;
            16'd16589: data <= 8'h07;
            16'd16590: data <= 8'hE0;
            16'd16591: data <= 8'h07;
            16'd16592: data <= 8'hE0;
            16'd16593: data <= 8'h07;
            16'd16594: data <= 8'hE0;
            16'd16595: data <= 8'h07;
            16'd16596: data <= 8'hE0;
            16'd16597: data <= 8'h07;
            16'd16598: data <= 8'hE0;
            16'd16599: data <= 8'h07;
            16'd16600: data <= 8'hFF;
            16'd16601: data <= 8'hFF;
            16'd16602: data <= 8'hE0;
            16'd16603: data <= 8'h07;
            16'd16604: data <= 8'hE0;
            16'd16605: data <= 8'h07;
            16'd16606: data <= 8'hE0;
            16'd16607: data <= 8'h07;
            16'd16608: data <= 8'hE0;
            16'd16609: data <= 8'h07;
            16'd16610: data <= 8'hE0;
            16'd16611: data <= 8'h07;
            16'd16612: data <= 8'hE0;
            16'd16613: data <= 8'h07;
            16'd16614: data <= 8'hE0;
            16'd16615: data <= 8'h07;
            16'd16616: data <= 8'hE0;
            16'd16617: data <= 8'h07;
            16'd16618: data <= 8'hE0;
            16'd16619: data <= 8'h07;
            16'd16620: data <= 8'hE0;
            16'd16621: data <= 8'h07;
            16'd16622: data <= 8'hE0;
            16'd16623: data <= 8'h07;
            16'd16624: data <= 8'hE0;
            16'd16625: data <= 8'h07;
            16'd16626: data <= 8'hE0;
            16'd16627: data <= 8'h07;
            16'd16628: data <= 8'hE0;
            16'd16629: data <= 8'h07;
            16'd16630: data <= 8'hE0;
            16'd16631: data <= 8'h07;
            16'd16632: data <= 8'hE0;
            16'd16633: data <= 8'h07;
            16'd16634: data <= 8'hE0;
            16'd16635: data <= 8'h07;
            16'd16636: data <= 8'hE0;
            16'd16637: data <= 8'h07;
            16'd16638: data <= 8'hE0;
            16'd16639: data <= 8'h07;
            16'd16640: data <= 8'hFF;
            16'd16641: data <= 8'hFF;
            16'd16642: data <= 8'hE0;
            16'd16643: data <= 8'h07;
            16'd16644: data <= 8'hE0;
            16'd16645: data <= 8'h07;
            16'd16646: data <= 8'hE0;
            16'd16647: data <= 8'h07;
            16'd16648: data <= 8'hE0;
            16'd16649: data <= 8'h07;
            16'd16650: data <= 8'hE0;
            16'd16651: data <= 8'h07;
            16'd16652: data <= 8'hE0;
            16'd16653: data <= 8'h07;
            16'd16654: data <= 8'hE0;
            16'd16655: data <= 8'h07;
            16'd16656: data <= 8'hE0;
            16'd16657: data <= 8'h07;
            16'd16658: data <= 8'hE0;
            16'd16659: data <= 8'h07;
            16'd16660: data <= 8'hE0;
            16'd16661: data <= 8'h07;
            16'd16662: data <= 8'hE0;
            16'd16663: data <= 8'h07;
            16'd16664: data <= 8'hE0;
            16'd16665: data <= 8'h07;
            16'd16666: data <= 8'hE0;
            16'd16667: data <= 8'h07;
            16'd16668: data <= 8'hE0;
            16'd16669: data <= 8'h07;
            16'd16670: data <= 8'hE0;
            16'd16671: data <= 8'h07;
            16'd16672: data <= 8'hE0;
            16'd16673: data <= 8'h07;
            16'd16674: data <= 8'hE0;
            16'd16675: data <= 8'h07;
            16'd16676: data <= 8'hE0;
            16'd16677: data <= 8'h07;
            16'd16678: data <= 8'hE0;
            16'd16679: data <= 8'h07;
            16'd16680: data <= 8'hFF;
            16'd16681: data <= 8'hFF;
            16'd16682: data <= 8'hE0;
            16'd16683: data <= 8'h07;
            16'd16684: data <= 8'hE0;
            16'd16685: data <= 8'h07;
            16'd16686: data <= 8'hE0;
            16'd16687: data <= 8'h07;
            16'd16688: data <= 8'hE0;
            16'd16689: data <= 8'h07;
            16'd16690: data <= 8'hE0;
            16'd16691: data <= 8'h07;
            16'd16692: data <= 8'hE0;
            16'd16693: data <= 8'h07;
            16'd16694: data <= 8'hE0;
            16'd16695: data <= 8'h07;
            16'd16696: data <= 8'hE0;
            16'd16697: data <= 8'h07;
            16'd16698: data <= 8'hE0;
            16'd16699: data <= 8'h07;
            16'd16700: data <= 8'hE0;
            16'd16701: data <= 8'h07;
            16'd16702: data <= 8'hE0;
            16'd16703: data <= 8'h07;
            16'd16704: data <= 8'hE0;
            16'd16705: data <= 8'h07;
            16'd16706: data <= 8'hE0;
            16'd16707: data <= 8'h07;
            16'd16708: data <= 8'hE0;
            16'd16709: data <= 8'h07;
            16'd16710: data <= 8'hE0;
            16'd16711: data <= 8'h07;
            16'd16712: data <= 8'hE0;
            16'd16713: data <= 8'h07;
            16'd16714: data <= 8'hE0;
            16'd16715: data <= 8'h07;
            16'd16716: data <= 8'hE0;
            16'd16717: data <= 8'h07;
            16'd16718: data <= 8'hE0;
            16'd16719: data <= 8'h07;
            16'd16720: data <= 8'hFF;
            16'd16721: data <= 8'hFF;
            16'd16722: data <= 8'hE0;
            16'd16723: data <= 8'h07;
            16'd16724: data <= 8'hE0;
            16'd16725: data <= 8'h07;
            16'd16726: data <= 8'hE0;
            16'd16727: data <= 8'h07;
            16'd16728: data <= 8'hE0;
            16'd16729: data <= 8'h07;
            16'd16730: data <= 8'hE0;
            16'd16731: data <= 8'h07;
            16'd16732: data <= 8'hE0;
            16'd16733: data <= 8'h07;
            16'd16734: data <= 8'hE0;
            16'd16735: data <= 8'h07;
            16'd16736: data <= 8'hE0;
            16'd16737: data <= 8'h07;
            16'd16738: data <= 8'hE0;
            16'd16739: data <= 8'h07;
            16'd16740: data <= 8'hE0;
            16'd16741: data <= 8'h07;
            16'd16742: data <= 8'hE0;
            16'd16743: data <= 8'h07;
            16'd16744: data <= 8'hE0;
            16'd16745: data <= 8'h07;
            16'd16746: data <= 8'hE0;
            16'd16747: data <= 8'h07;
            16'd16748: data <= 8'hE0;
            16'd16749: data <= 8'h07;
            16'd16750: data <= 8'hE0;
            16'd16751: data <= 8'h07;
            16'd16752: data <= 8'hE0;
            16'd16753: data <= 8'h07;
            16'd16754: data <= 8'hE0;
            16'd16755: data <= 8'h07;
            16'd16756: data <= 8'hE0;
            16'd16757: data <= 8'h07;
            16'd16758: data <= 8'hE0;
            16'd16759: data <= 8'h07;
            16'd16760: data <= 8'hFF;
            16'd16761: data <= 8'hFF;
            16'd16762: data <= 8'hE0;
            16'd16763: data <= 8'h07;
            16'd16764: data <= 8'hE0;
            16'd16765: data <= 8'h07;
            16'd16766: data <= 8'hE0;
            16'd16767: data <= 8'h07;
            16'd16768: data <= 8'hE0;
            16'd16769: data <= 8'h07;
            16'd16770: data <= 8'hE0;
            16'd16771: data <= 8'h07;
            16'd16772: data <= 8'hE0;
            16'd16773: data <= 8'h07;
            16'd16774: data <= 8'hE0;
            16'd16775: data <= 8'h07;
            16'd16776: data <= 8'hE0;
            16'd16777: data <= 8'h07;
            16'd16778: data <= 8'hE0;
            16'd16779: data <= 8'h07;
            16'd16780: data <= 8'hE0;
            16'd16781: data <= 8'h07;
            16'd16782: data <= 8'hE0;
            16'd16783: data <= 8'h07;
            16'd16784: data <= 8'hE0;
            16'd16785: data <= 8'h07;
            16'd16786: data <= 8'hE0;
            16'd16787: data <= 8'h07;
            16'd16788: data <= 8'hE0;
            16'd16789: data <= 8'h07;
            16'd16790: data <= 8'hE0;
            16'd16791: data <= 8'h07;
            16'd16792: data <= 8'hE0;
            16'd16793: data <= 8'h07;
            16'd16794: data <= 8'hE0;
            16'd16795: data <= 8'h07;
            16'd16796: data <= 8'hE0;
            16'd16797: data <= 8'h07;
            16'd16798: data <= 8'hE0;
            16'd16799: data <= 8'h07;
            16'd16800: data <= 8'hFF;
            16'd16801: data <= 8'hFF;
            16'd16802: data <= 8'hE0;
            16'd16803: data <= 8'h07;
            16'd16804: data <= 8'hE0;
            16'd16805: data <= 8'h07;
            16'd16806: data <= 8'hE0;
            16'd16807: data <= 8'h07;
            16'd16808: data <= 8'hE0;
            16'd16809: data <= 8'h07;
            16'd16810: data <= 8'hE0;
            16'd16811: data <= 8'h07;
            16'd16812: data <= 8'hE0;
            16'd16813: data <= 8'h07;
            16'd16814: data <= 8'hE0;
            16'd16815: data <= 8'h07;
            16'd16816: data <= 8'hE0;
            16'd16817: data <= 8'h07;
            16'd16818: data <= 8'hE0;
            16'd16819: data <= 8'h07;
            16'd16820: data <= 8'hE0;
            16'd16821: data <= 8'h07;
            16'd16822: data <= 8'hE0;
            16'd16823: data <= 8'h07;
            16'd16824: data <= 8'hE0;
            16'd16825: data <= 8'h07;
            16'd16826: data <= 8'hE0;
            16'd16827: data <= 8'h07;
            16'd16828: data <= 8'hE0;
            16'd16829: data <= 8'h07;
            16'd16830: data <= 8'hE0;
            16'd16831: data <= 8'h07;
            16'd16832: data <= 8'hE0;
            16'd16833: data <= 8'h07;
            16'd16834: data <= 8'hE0;
            16'd16835: data <= 8'h07;
            16'd16836: data <= 8'hE0;
            16'd16837: data <= 8'h07;
            16'd16838: data <= 8'hE0;
            16'd16839: data <= 8'h07;
            16'd16840: data <= 8'hFF;
            16'd16841: data <= 8'hFF;
            16'd16842: data <= 8'hE0;
            16'd16843: data <= 8'h07;
            16'd16844: data <= 8'hE0;
            16'd16845: data <= 8'h07;
            16'd16846: data <= 8'hE0;
            16'd16847: data <= 8'h07;
            16'd16848: data <= 8'hE0;
            16'd16849: data <= 8'h07;
            16'd16850: data <= 8'hE0;
            16'd16851: data <= 8'h07;
            16'd16852: data <= 8'hE0;
            16'd16853: data <= 8'h07;
            16'd16854: data <= 8'hE0;
            16'd16855: data <= 8'h07;
            16'd16856: data <= 8'hE0;
            16'd16857: data <= 8'h07;
            16'd16858: data <= 8'hE0;
            16'd16859: data <= 8'h07;
            16'd16860: data <= 8'hE0;
            16'd16861: data <= 8'h07;
            16'd16862: data <= 8'hE0;
            16'd16863: data <= 8'h07;
            16'd16864: data <= 8'hE0;
            16'd16865: data <= 8'h07;
            16'd16866: data <= 8'hE0;
            16'd16867: data <= 8'h07;
            16'd16868: data <= 8'hE0;
            16'd16869: data <= 8'h07;
            16'd16870: data <= 8'hE0;
            16'd16871: data <= 8'h07;
            16'd16872: data <= 8'hE0;
            16'd16873: data <= 8'h07;
            16'd16874: data <= 8'hE0;
            16'd16875: data <= 8'h07;
            16'd16876: data <= 8'hE0;
            16'd16877: data <= 8'h07;
            16'd16878: data <= 8'hE0;
            16'd16879: data <= 8'h07;
            16'd16880: data <= 8'hFF;
            16'd16881: data <= 8'hFF;
            16'd16882: data <= 8'hE0;
            16'd16883: data <= 8'h07;
            16'd16884: data <= 8'hE0;
            16'd16885: data <= 8'h07;
            16'd16886: data <= 8'hE0;
            16'd16887: data <= 8'h07;
            16'd16888: data <= 8'hE0;
            16'd16889: data <= 8'h07;
            16'd16890: data <= 8'hE0;
            16'd16891: data <= 8'h07;
            16'd16892: data <= 8'hE0;
            16'd16893: data <= 8'h07;
            16'd16894: data <= 8'hE0;
            16'd16895: data <= 8'h07;
            16'd16896: data <= 8'hE0;
            16'd16897: data <= 8'h07;
            16'd16898: data <= 8'hE0;
            16'd16899: data <= 8'h07;
            16'd16900: data <= 8'hE0;
            16'd16901: data <= 8'h07;
            16'd16902: data <= 8'hE0;
            16'd16903: data <= 8'h07;
            16'd16904: data <= 8'hE0;
            16'd16905: data <= 8'h07;
            16'd16906: data <= 8'hE0;
            16'd16907: data <= 8'h07;
            16'd16908: data <= 8'hE0;
            16'd16909: data <= 8'h07;
            16'd16910: data <= 8'hE0;
            16'd16911: data <= 8'h07;
            16'd16912: data <= 8'hE0;
            16'd16913: data <= 8'h07;
            16'd16914: data <= 8'hE0;
            16'd16915: data <= 8'h07;
            16'd16916: data <= 8'hE0;
            16'd16917: data <= 8'h07;
            16'd16918: data <= 8'hE0;
            16'd16919: data <= 8'h07;
            16'd16920: data <= 8'hFF;
            16'd16921: data <= 8'hFF;
            16'd16922: data <= 8'hE0;
            16'd16923: data <= 8'h07;
            16'd16924: data <= 8'hE0;
            16'd16925: data <= 8'h07;
            16'd16926: data <= 8'hE0;
            16'd16927: data <= 8'h07;
            16'd16928: data <= 8'hE0;
            16'd16929: data <= 8'h07;
            16'd16930: data <= 8'hE0;
            16'd16931: data <= 8'h07;
            16'd16932: data <= 8'hE0;
            16'd16933: data <= 8'h07;
            16'd16934: data <= 8'hE0;
            16'd16935: data <= 8'h07;
            16'd16936: data <= 8'hE0;
            16'd16937: data <= 8'h07;
            16'd16938: data <= 8'hE0;
            16'd16939: data <= 8'h07;
            16'd16940: data <= 8'hE0;
            16'd16941: data <= 8'h07;
            16'd16942: data <= 8'hE0;
            16'd16943: data <= 8'h07;
            16'd16944: data <= 8'hE0;
            16'd16945: data <= 8'h07;
            16'd16946: data <= 8'hE0;
            16'd16947: data <= 8'h07;
            16'd16948: data <= 8'hE0;
            16'd16949: data <= 8'h07;
            16'd16950: data <= 8'hE0;
            16'd16951: data <= 8'h07;
            16'd16952: data <= 8'hE0;
            16'd16953: data <= 8'h07;
            16'd16954: data <= 8'hE0;
            16'd16955: data <= 8'h07;
            16'd16956: data <= 8'hE0;
            16'd16957: data <= 8'h07;
            16'd16958: data <= 8'hE0;
            16'd16959: data <= 8'h07;
            16'd16960: data <= 8'hFF;
            16'd16961: data <= 8'hFF;
            16'd16962: data <= 8'hE0;
            16'd16963: data <= 8'h07;
            16'd16964: data <= 8'hE0;
            16'd16965: data <= 8'h07;
            16'd16966: data <= 8'hE0;
            16'd16967: data <= 8'h07;
            16'd16968: data <= 8'hE0;
            16'd16969: data <= 8'h07;
            16'd16970: data <= 8'hE0;
            16'd16971: data <= 8'h07;
            16'd16972: data <= 8'hE0;
            16'd16973: data <= 8'h07;
            16'd16974: data <= 8'hE0;
            16'd16975: data <= 8'h07;
            16'd16976: data <= 8'hE0;
            16'd16977: data <= 8'h07;
            16'd16978: data <= 8'hE0;
            16'd16979: data <= 8'h07;
            16'd16980: data <= 8'hE0;
            16'd16981: data <= 8'h07;
            16'd16982: data <= 8'hE0;
            16'd16983: data <= 8'h07;
            16'd16984: data <= 8'hE0;
            16'd16985: data <= 8'h07;
            16'd16986: data <= 8'hE0;
            16'd16987: data <= 8'h07;
            16'd16988: data <= 8'hE0;
            16'd16989: data <= 8'h07;
            16'd16990: data <= 8'hE0;
            16'd16991: data <= 8'h07;
            16'd16992: data <= 8'hE0;
            16'd16993: data <= 8'h07;
            16'd16994: data <= 8'hE0;
            16'd16995: data <= 8'h07;
            16'd16996: data <= 8'hE0;
            16'd16997: data <= 8'h07;
            16'd16998: data <= 8'hE0;
            16'd16999: data <= 8'h07;
            16'd17000: data <= 8'hFF;
            16'd17001: data <= 8'hFF;
            16'd17002: data <= 8'hE0;
            16'd17003: data <= 8'h07;
            16'd17004: data <= 8'hE0;
            16'd17005: data <= 8'h07;
            16'd17006: data <= 8'hE0;
            16'd17007: data <= 8'h07;
            16'd17008: data <= 8'hE0;
            16'd17009: data <= 8'h07;
            16'd17010: data <= 8'hE0;
            16'd17011: data <= 8'h07;
            16'd17012: data <= 8'hE0;
            16'd17013: data <= 8'h07;
            16'd17014: data <= 8'hE0;
            16'd17015: data <= 8'h07;
            16'd17016: data <= 8'hE0;
            16'd17017: data <= 8'h07;
            16'd17018: data <= 8'hE0;
            16'd17019: data <= 8'h07;
            16'd17020: data <= 8'hE0;
            16'd17021: data <= 8'h07;
            16'd17022: data <= 8'hE0;
            16'd17023: data <= 8'h07;
            16'd17024: data <= 8'hE0;
            16'd17025: data <= 8'h07;
            16'd17026: data <= 8'hE0;
            16'd17027: data <= 8'h07;
            16'd17028: data <= 8'hE0;
            16'd17029: data <= 8'h07;
            16'd17030: data <= 8'hE0;
            16'd17031: data <= 8'h07;
            16'd17032: data <= 8'hE0;
            16'd17033: data <= 8'h07;
            16'd17034: data <= 8'hE0;
            16'd17035: data <= 8'h07;
            16'd17036: data <= 8'hE0;
            16'd17037: data <= 8'h07;
            16'd17038: data <= 8'hE0;
            16'd17039: data <= 8'h07;
            16'd17040: data <= 8'hFF;
            16'd17041: data <= 8'hFF;
            16'd17042: data <= 8'hE0;
            16'd17043: data <= 8'h07;
            16'd17044: data <= 8'hE0;
            16'd17045: data <= 8'h07;
            16'd17046: data <= 8'hE0;
            16'd17047: data <= 8'h07;
            16'd17048: data <= 8'hE0;
            16'd17049: data <= 8'h07;
            16'd17050: data <= 8'hE0;
            16'd17051: data <= 8'h07;
            16'd17052: data <= 8'hE0;
            16'd17053: data <= 8'h07;
            16'd17054: data <= 8'hE0;
            16'd17055: data <= 8'h07;
            16'd17056: data <= 8'hE0;
            16'd17057: data <= 8'h07;
            16'd17058: data <= 8'hE0;
            16'd17059: data <= 8'h07;
            16'd17060: data <= 8'hE0;
            16'd17061: data <= 8'h07;
            16'd17062: data <= 8'hE0;
            16'd17063: data <= 8'h07;
            16'd17064: data <= 8'hE0;
            16'd17065: data <= 8'h07;
            16'd17066: data <= 8'hE0;
            16'd17067: data <= 8'h07;
            16'd17068: data <= 8'hE0;
            16'd17069: data <= 8'h07;
            16'd17070: data <= 8'hE0;
            16'd17071: data <= 8'h07;
            16'd17072: data <= 8'hE0;
            16'd17073: data <= 8'h07;
            16'd17074: data <= 8'hE0;
            16'd17075: data <= 8'h07;
            16'd17076: data <= 8'hE0;
            16'd17077: data <= 8'h07;
            16'd17078: data <= 8'hE0;
            16'd17079: data <= 8'h07;
            16'd17080: data <= 8'hFF;
            16'd17081: data <= 8'hFF;
            16'd17082: data <= 8'hE0;
            16'd17083: data <= 8'h07;
            16'd17084: data <= 8'hE0;
            16'd17085: data <= 8'h07;
            16'd17086: data <= 8'hE0;
            16'd17087: data <= 8'h07;
            16'd17088: data <= 8'hE0;
            16'd17089: data <= 8'h07;
            16'd17090: data <= 8'hE0;
            16'd17091: data <= 8'h07;
            16'd17092: data <= 8'hE0;
            16'd17093: data <= 8'h07;
            16'd17094: data <= 8'hE0;
            16'd17095: data <= 8'h07;
            16'd17096: data <= 8'hE0;
            16'd17097: data <= 8'h07;
            16'd17098: data <= 8'hE0;
            16'd17099: data <= 8'h07;
            16'd17100: data <= 8'hE0;
            16'd17101: data <= 8'h07;
            16'd17102: data <= 8'hE0;
            16'd17103: data <= 8'h07;
            16'd17104: data <= 8'hE0;
            16'd17105: data <= 8'h07;
            16'd17106: data <= 8'hE0;
            16'd17107: data <= 8'h07;
            16'd17108: data <= 8'hE0;
            16'd17109: data <= 8'h07;
            16'd17110: data <= 8'hE0;
            16'd17111: data <= 8'h07;
            16'd17112: data <= 8'hE0;
            16'd17113: data <= 8'h07;
            16'd17114: data <= 8'hE0;
            16'd17115: data <= 8'h07;
            16'd17116: data <= 8'hE0;
            16'd17117: data <= 8'h07;
            16'd17118: data <= 8'hE0;
            16'd17119: data <= 8'h07;
            16'd17120: data <= 8'hFF;
            16'd17121: data <= 8'hFF;
            16'd17122: data <= 8'hE0;
            16'd17123: data <= 8'h07;
            16'd17124: data <= 8'hE0;
            16'd17125: data <= 8'h07;
            16'd17126: data <= 8'hE0;
            16'd17127: data <= 8'h07;
            16'd17128: data <= 8'hE0;
            16'd17129: data <= 8'h07;
            16'd17130: data <= 8'hE0;
            16'd17131: data <= 8'h07;
            16'd17132: data <= 8'hE0;
            16'd17133: data <= 8'h07;
            16'd17134: data <= 8'hE0;
            16'd17135: data <= 8'h07;
            16'd17136: data <= 8'hE0;
            16'd17137: data <= 8'h07;
            16'd17138: data <= 8'hE0;
            16'd17139: data <= 8'h07;
            16'd17140: data <= 8'hE0;
            16'd17141: data <= 8'h07;
            16'd17142: data <= 8'hE0;
            16'd17143: data <= 8'h07;
            16'd17144: data <= 8'hE0;
            16'd17145: data <= 8'h07;
            16'd17146: data <= 8'hE0;
            16'd17147: data <= 8'h07;
            16'd17148: data <= 8'hE0;
            16'd17149: data <= 8'h07;
            16'd17150: data <= 8'hE0;
            16'd17151: data <= 8'h07;
            16'd17152: data <= 8'hE0;
            16'd17153: data <= 8'h07;
            16'd17154: data <= 8'hE0;
            16'd17155: data <= 8'h07;
            16'd17156: data <= 8'hE0;
            16'd17157: data <= 8'h07;
            16'd17158: data <= 8'hE0;
            16'd17159: data <= 8'h07;
            16'd17160: data <= 8'hFF;
            16'd17161: data <= 8'hFF;
            16'd17162: data <= 8'hE0;
            16'd17163: data <= 8'h07;
            16'd17164: data <= 8'hE0;
            16'd17165: data <= 8'h07;
            16'd17166: data <= 8'hE0;
            16'd17167: data <= 8'h07;
            16'd17168: data <= 8'hE0;
            16'd17169: data <= 8'h07;
            16'd17170: data <= 8'hE0;
            16'd17171: data <= 8'h07;
            16'd17172: data <= 8'hE0;
            16'd17173: data <= 8'h07;
            16'd17174: data <= 8'hE0;
            16'd17175: data <= 8'h07;
            16'd17176: data <= 8'hE0;
            16'd17177: data <= 8'h07;
            16'd17178: data <= 8'hE0;
            16'd17179: data <= 8'h07;
            16'd17180: data <= 8'hE0;
            16'd17181: data <= 8'h07;
            16'd17182: data <= 8'hE0;
            16'd17183: data <= 8'h07;
            16'd17184: data <= 8'hE0;
            16'd17185: data <= 8'h07;
            16'd17186: data <= 8'hE0;
            16'd17187: data <= 8'h07;
            16'd17188: data <= 8'hE0;
            16'd17189: data <= 8'h07;
            16'd17190: data <= 8'hE0;
            16'd17191: data <= 8'h07;
            16'd17192: data <= 8'hE0;
            16'd17193: data <= 8'h07;
            16'd17194: data <= 8'hE0;
            16'd17195: data <= 8'h07;
            16'd17196: data <= 8'hE0;
            16'd17197: data <= 8'h07;
            16'd17198: data <= 8'hE0;
            16'd17199: data <= 8'h07;
            16'd17200: data <= 8'hFF;
            16'd17201: data <= 8'hFF;
            16'd17202: data <= 8'hE0;
            16'd17203: data <= 8'h07;
            16'd17204: data <= 8'hE0;
            16'd17205: data <= 8'h07;
            16'd17206: data <= 8'hE0;
            16'd17207: data <= 8'h07;
            16'd17208: data <= 8'hE0;
            16'd17209: data <= 8'h07;
            16'd17210: data <= 8'hE0;
            16'd17211: data <= 8'h07;
            16'd17212: data <= 8'hE0;
            16'd17213: data <= 8'h07;
            16'd17214: data <= 8'hE0;
            16'd17215: data <= 8'h07;
            16'd17216: data <= 8'hE0;
            16'd17217: data <= 8'h07;
            16'd17218: data <= 8'hE0;
            16'd17219: data <= 8'h07;
            16'd17220: data <= 8'hE0;
            16'd17221: data <= 8'h07;
            16'd17222: data <= 8'hE0;
            16'd17223: data <= 8'h07;
            16'd17224: data <= 8'hE0;
            16'd17225: data <= 8'h07;
            16'd17226: data <= 8'hE0;
            16'd17227: data <= 8'h07;
            16'd17228: data <= 8'hE0;
            16'd17229: data <= 8'h07;
            16'd17230: data <= 8'hE0;
            16'd17231: data <= 8'h07;
            16'd17232: data <= 8'hE0;
            16'd17233: data <= 8'h07;
            16'd17234: data <= 8'hE0;
            16'd17235: data <= 8'h07;
            16'd17236: data <= 8'hE0;
            16'd17237: data <= 8'h07;
            16'd17238: data <= 8'hE0;
            16'd17239: data <= 8'h07;
            16'd17240: data <= 8'hFF;
            16'd17241: data <= 8'hFF;
            16'd17242: data <= 8'hE0;
            16'd17243: data <= 8'h07;
            16'd17244: data <= 8'hE0;
            16'd17245: data <= 8'h07;
            16'd17246: data <= 8'hE0;
            16'd17247: data <= 8'h07;
            16'd17248: data <= 8'hE0;
            16'd17249: data <= 8'h07;
            16'd17250: data <= 8'hE0;
            16'd17251: data <= 8'h07;
            16'd17252: data <= 8'hE0;
            16'd17253: data <= 8'h07;
            16'd17254: data <= 8'hE0;
            16'd17255: data <= 8'h07;
            16'd17256: data <= 8'hE0;
            16'd17257: data <= 8'h07;
            16'd17258: data <= 8'hE0;
            16'd17259: data <= 8'h07;
            16'd17260: data <= 8'hE0;
            16'd17261: data <= 8'h07;
            16'd17262: data <= 8'hE0;
            16'd17263: data <= 8'h07;
            16'd17264: data <= 8'hE0;
            16'd17265: data <= 8'h07;
            16'd17266: data <= 8'hE0;
            16'd17267: data <= 8'h07;
            16'd17268: data <= 8'hE0;
            16'd17269: data <= 8'h07;
            16'd17270: data <= 8'hE0;
            16'd17271: data <= 8'h07;
            16'd17272: data <= 8'hE0;
            16'd17273: data <= 8'h07;
            16'd17274: data <= 8'hE0;
            16'd17275: data <= 8'h07;
            16'd17276: data <= 8'hE0;
            16'd17277: data <= 8'h07;
            16'd17278: data <= 8'hE0;
            16'd17279: data <= 8'h07;
            16'd17280: data <= 8'hFF;
            16'd17281: data <= 8'hFF;
            16'd17282: data <= 8'hE0;
            16'd17283: data <= 8'h07;
            16'd17284: data <= 8'hE0;
            16'd17285: data <= 8'h07;
            16'd17286: data <= 8'hE0;
            16'd17287: data <= 8'h07;
            16'd17288: data <= 8'hE0;
            16'd17289: data <= 8'h07;
            16'd17290: data <= 8'hE0;
            16'd17291: data <= 8'h07;
            16'd17292: data <= 8'hE0;
            16'd17293: data <= 8'h07;
            16'd17294: data <= 8'hE0;
            16'd17295: data <= 8'h07;
            16'd17296: data <= 8'hE0;
            16'd17297: data <= 8'h07;
            16'd17298: data <= 8'hE0;
            16'd17299: data <= 8'h07;
            16'd17300: data <= 8'hE0;
            16'd17301: data <= 8'h07;
            16'd17302: data <= 8'hE0;
            16'd17303: data <= 8'h07;
            16'd17304: data <= 8'hE0;
            16'd17305: data <= 8'h07;
            16'd17306: data <= 8'hE0;
            16'd17307: data <= 8'h07;
            16'd17308: data <= 8'hE0;
            16'd17309: data <= 8'h07;
            16'd17310: data <= 8'hE0;
            16'd17311: data <= 8'h07;
            16'd17312: data <= 8'hE0;
            16'd17313: data <= 8'h07;
            16'd17314: data <= 8'hE0;
            16'd17315: data <= 8'h07;
            16'd17316: data <= 8'hE0;
            16'd17317: data <= 8'h07;
            16'd17318: data <= 8'hE0;
            16'd17319: data <= 8'h07;
            16'd17320: data <= 8'hFF;
            16'd17321: data <= 8'hFF;
            16'd17322: data <= 8'hE0;
            16'd17323: data <= 8'h07;
            16'd17324: data <= 8'hE0;
            16'd17325: data <= 8'h07;
            16'd17326: data <= 8'hE0;
            16'd17327: data <= 8'h07;
            16'd17328: data <= 8'hE0;
            16'd17329: data <= 8'h07;
            16'd17330: data <= 8'hE0;
            16'd17331: data <= 8'h07;
            16'd17332: data <= 8'hE0;
            16'd17333: data <= 8'h07;
            16'd17334: data <= 8'hE0;
            16'd17335: data <= 8'h07;
            16'd17336: data <= 8'hE0;
            16'd17337: data <= 8'h07;
            16'd17338: data <= 8'hE0;
            16'd17339: data <= 8'h07;
            16'd17340: data <= 8'hE0;
            16'd17341: data <= 8'h07;
            16'd17342: data <= 8'hE0;
            16'd17343: data <= 8'h07;
            16'd17344: data <= 8'hE0;
            16'd17345: data <= 8'h07;
            16'd17346: data <= 8'hE0;
            16'd17347: data <= 8'h07;
            16'd17348: data <= 8'hE0;
            16'd17349: data <= 8'h07;
            16'd17350: data <= 8'hE0;
            16'd17351: data <= 8'h07;
            16'd17352: data <= 8'hE0;
            16'd17353: data <= 8'h07;
            16'd17354: data <= 8'hE0;
            16'd17355: data <= 8'h07;
            16'd17356: data <= 8'hE0;
            16'd17357: data <= 8'h07;
            16'd17358: data <= 8'hE0;
            16'd17359: data <= 8'h07;
            16'd17360: data <= 8'hFF;
            16'd17361: data <= 8'hFF;
            16'd17362: data <= 8'hE0;
            16'd17363: data <= 8'h07;
            16'd17364: data <= 8'hE0;
            16'd17365: data <= 8'h07;
            16'd17366: data <= 8'hE0;
            16'd17367: data <= 8'h07;
            16'd17368: data <= 8'hE0;
            16'd17369: data <= 8'h07;
            16'd17370: data <= 8'hE0;
            16'd17371: data <= 8'h07;
            16'd17372: data <= 8'hE0;
            16'd17373: data <= 8'h07;
            16'd17374: data <= 8'hE0;
            16'd17375: data <= 8'h07;
            16'd17376: data <= 8'hE0;
            16'd17377: data <= 8'h07;
            16'd17378: data <= 8'hE0;
            16'd17379: data <= 8'h07;
            16'd17380: data <= 8'hE0;
            16'd17381: data <= 8'h07;
            16'd17382: data <= 8'hE0;
            16'd17383: data <= 8'h07;
            16'd17384: data <= 8'hE0;
            16'd17385: data <= 8'h07;
            16'd17386: data <= 8'hE0;
            16'd17387: data <= 8'h07;
            16'd17388: data <= 8'hE0;
            16'd17389: data <= 8'h07;
            16'd17390: data <= 8'hE0;
            16'd17391: data <= 8'h07;
            16'd17392: data <= 8'hE0;
            16'd17393: data <= 8'h07;
            16'd17394: data <= 8'hE0;
            16'd17395: data <= 8'h07;
            16'd17396: data <= 8'hE0;
            16'd17397: data <= 8'h07;
            16'd17398: data <= 8'hE0;
            16'd17399: data <= 8'h07;
            16'd17400: data <= 8'hFF;
            16'd17401: data <= 8'hFF;
            16'd17402: data <= 8'hE0;
            16'd17403: data <= 8'h07;
            16'd17404: data <= 8'hE0;
            16'd17405: data <= 8'h07;
            16'd17406: data <= 8'hE0;
            16'd17407: data <= 8'h07;
            16'd17408: data <= 8'hE0;
            16'd17409: data <= 8'h07;
            16'd17410: data <= 8'hE0;
            16'd17411: data <= 8'h07;
            16'd17412: data <= 8'hE0;
            16'd17413: data <= 8'h07;
            16'd17414: data <= 8'hE0;
            16'd17415: data <= 8'h07;
            16'd17416: data <= 8'hE0;
            16'd17417: data <= 8'h07;
            16'd17418: data <= 8'hE0;
            16'd17419: data <= 8'h07;
            16'd17420: data <= 8'hE0;
            16'd17421: data <= 8'h07;
            16'd17422: data <= 8'hE0;
            16'd17423: data <= 8'h07;
            16'd17424: data <= 8'hE0;
            16'd17425: data <= 8'h07;
            16'd17426: data <= 8'hE0;
            16'd17427: data <= 8'h07;
            16'd17428: data <= 8'hE0;
            16'd17429: data <= 8'h07;
            16'd17430: data <= 8'hE0;
            16'd17431: data <= 8'h07;
            16'd17432: data <= 8'hE0;
            16'd17433: data <= 8'h07;
            16'd17434: data <= 8'hE0;
            16'd17435: data <= 8'h07;
            16'd17436: data <= 8'hE0;
            16'd17437: data <= 8'h07;
            16'd17438: data <= 8'hE0;
            16'd17439: data <= 8'h07;
            16'd17440: data <= 8'hFF;
            16'd17441: data <= 8'hFF;
            16'd17442: data <= 8'hE0;
            16'd17443: data <= 8'h07;
            16'd17444: data <= 8'hE0;
            16'd17445: data <= 8'h07;
            16'd17446: data <= 8'hE0;
            16'd17447: data <= 8'h07;
            16'd17448: data <= 8'hE0;
            16'd17449: data <= 8'h07;
            16'd17450: data <= 8'hE0;
            16'd17451: data <= 8'h07;
            16'd17452: data <= 8'hE0;
            16'd17453: data <= 8'h07;
            16'd17454: data <= 8'hE0;
            16'd17455: data <= 8'h07;
            16'd17456: data <= 8'hE0;
            16'd17457: data <= 8'h07;
            16'd17458: data <= 8'hE0;
            16'd17459: data <= 8'h07;
            16'd17460: data <= 8'hE0;
            16'd17461: data <= 8'h07;
            16'd17462: data <= 8'hE0;
            16'd17463: data <= 8'h07;
            16'd17464: data <= 8'hE0;
            16'd17465: data <= 8'h07;
            16'd17466: data <= 8'hE0;
            16'd17467: data <= 8'h07;
            16'd17468: data <= 8'hE0;
            16'd17469: data <= 8'h07;
            16'd17470: data <= 8'hE0;
            16'd17471: data <= 8'h07;
            16'd17472: data <= 8'hE0;
            16'd17473: data <= 8'h07;
            16'd17474: data <= 8'hE0;
            16'd17475: data <= 8'h07;
            16'd17476: data <= 8'hE0;
            16'd17477: data <= 8'h07;
            16'd17478: data <= 8'hE0;
            16'd17479: data <= 8'h07;
            16'd17480: data <= 8'hFF;
            16'd17481: data <= 8'hFF;
            16'd17482: data <= 8'hE0;
            16'd17483: data <= 8'h07;
            16'd17484: data <= 8'hE0;
            16'd17485: data <= 8'h07;
            16'd17486: data <= 8'hE0;
            16'd17487: data <= 8'h07;
            16'd17488: data <= 8'hE0;
            16'd17489: data <= 8'h07;
            16'd17490: data <= 8'hE0;
            16'd17491: data <= 8'h07;
            16'd17492: data <= 8'hE0;
            16'd17493: data <= 8'h07;
            16'd17494: data <= 8'hE0;
            16'd17495: data <= 8'h07;
            16'd17496: data <= 8'hE0;
            16'd17497: data <= 8'h07;
            16'd17498: data <= 8'hE0;
            16'd17499: data <= 8'h07;
            16'd17500: data <= 8'hE0;
            16'd17501: data <= 8'h07;
            16'd17502: data <= 8'hE0;
            16'd17503: data <= 8'h07;
            16'd17504: data <= 8'hE0;
            16'd17505: data <= 8'h07;
            16'd17506: data <= 8'hE0;
            16'd17507: data <= 8'h07;
            16'd17508: data <= 8'hE0;
            16'd17509: data <= 8'h07;
            16'd17510: data <= 8'hE0;
            16'd17511: data <= 8'h07;
            16'd17512: data <= 8'hE0;
            16'd17513: data <= 8'h07;
            16'd17514: data <= 8'hE0;
            16'd17515: data <= 8'h07;
            16'd17516: data <= 8'hE0;
            16'd17517: data <= 8'h07;
            16'd17518: data <= 8'hE0;
            16'd17519: data <= 8'h07;
            16'd17520: data <= 8'hFF;
            16'd17521: data <= 8'hFF;
            16'd17522: data <= 8'hE0;
            16'd17523: data <= 8'h07;
            16'd17524: data <= 8'hE0;
            16'd17525: data <= 8'h07;
            16'd17526: data <= 8'hE0;
            16'd17527: data <= 8'h07;
            16'd17528: data <= 8'hE0;
            16'd17529: data <= 8'h07;
            16'd17530: data <= 8'hE0;
            16'd17531: data <= 8'h07;
            16'd17532: data <= 8'hE0;
            16'd17533: data <= 8'h07;
            16'd17534: data <= 8'hE0;
            16'd17535: data <= 8'h07;
            16'd17536: data <= 8'hE0;
            16'd17537: data <= 8'h07;
            16'd17538: data <= 8'hE0;
            16'd17539: data <= 8'h07;
            16'd17540: data <= 8'hE0;
            16'd17541: data <= 8'h07;
            16'd17542: data <= 8'hE0;
            16'd17543: data <= 8'h07;
            16'd17544: data <= 8'hE0;
            16'd17545: data <= 8'h07;
            16'd17546: data <= 8'hE0;
            16'd17547: data <= 8'h07;
            16'd17548: data <= 8'hE0;
            16'd17549: data <= 8'h07;
            16'd17550: data <= 8'hE0;
            16'd17551: data <= 8'h07;
            16'd17552: data <= 8'hE0;
            16'd17553: data <= 8'h07;
            16'd17554: data <= 8'hE0;
            16'd17555: data <= 8'h07;
            16'd17556: data <= 8'hE0;
            16'd17557: data <= 8'h07;
            16'd17558: data <= 8'hE0;
            16'd17559: data <= 8'h07;
            16'd17560: data <= 8'hFF;
            16'd17561: data <= 8'hFF;
            16'd17562: data <= 8'hE0;
            16'd17563: data <= 8'h07;
            16'd17564: data <= 8'hE0;
            16'd17565: data <= 8'h07;
            16'd17566: data <= 8'hE0;
            16'd17567: data <= 8'h07;
            16'd17568: data <= 8'hE0;
            16'd17569: data <= 8'h07;
            16'd17570: data <= 8'hE0;
            16'd17571: data <= 8'h07;
            16'd17572: data <= 8'hE0;
            16'd17573: data <= 8'h07;
            16'd17574: data <= 8'hE0;
            16'd17575: data <= 8'h07;
            16'd17576: data <= 8'hE0;
            16'd17577: data <= 8'h07;
            16'd17578: data <= 8'hE0;
            16'd17579: data <= 8'h07;
            16'd17580: data <= 8'hE0;
            16'd17581: data <= 8'h07;
            16'd17582: data <= 8'hE0;
            16'd17583: data <= 8'h07;
            16'd17584: data <= 8'hE0;
            16'd17585: data <= 8'h07;
            16'd17586: data <= 8'hE0;
            16'd17587: data <= 8'h07;
            16'd17588: data <= 8'hE0;
            16'd17589: data <= 8'h07;
            16'd17590: data <= 8'hE0;
            16'd17591: data <= 8'h07;
            16'd17592: data <= 8'hE0;
            16'd17593: data <= 8'h07;
            16'd17594: data <= 8'hE0;
            16'd17595: data <= 8'h07;
            16'd17596: data <= 8'hE0;
            16'd17597: data <= 8'h07;
            16'd17598: data <= 8'hE0;
            16'd17599: data <= 8'h07;
            16'd17600: data <= 8'hFF;
            16'd17601: data <= 8'hFF;
            16'd17602: data <= 8'hE0;
            16'd17603: data <= 8'h07;
            16'd17604: data <= 8'hE0;
            16'd17605: data <= 8'h07;
            16'd17606: data <= 8'hE0;
            16'd17607: data <= 8'h07;
            16'd17608: data <= 8'hE0;
            16'd17609: data <= 8'h07;
            16'd17610: data <= 8'hE0;
            16'd17611: data <= 8'h07;
            16'd17612: data <= 8'hE0;
            16'd17613: data <= 8'h07;
            16'd17614: data <= 8'hE0;
            16'd17615: data <= 8'h07;
            16'd17616: data <= 8'hE0;
            16'd17617: data <= 8'h07;
            16'd17618: data <= 8'hE0;
            16'd17619: data <= 8'h07;
            16'd17620: data <= 8'hE0;
            16'd17621: data <= 8'h07;
            16'd17622: data <= 8'hE0;
            16'd17623: data <= 8'h07;
            16'd17624: data <= 8'hE0;
            16'd17625: data <= 8'h07;
            16'd17626: data <= 8'hE0;
            16'd17627: data <= 8'h07;
            16'd17628: data <= 8'hE0;
            16'd17629: data <= 8'h07;
            16'd17630: data <= 8'hE0;
            16'd17631: data <= 8'h07;
            16'd17632: data <= 8'hE0;
            16'd17633: data <= 8'h07;
            16'd17634: data <= 8'hE0;
            16'd17635: data <= 8'h07;
            16'd17636: data <= 8'hE0;
            16'd17637: data <= 8'h07;
            16'd17638: data <= 8'hE0;
            16'd17639: data <= 8'h07;
            16'd17640: data <= 8'hFF;
            16'd17641: data <= 8'hFF;
            16'd17642: data <= 8'hE0;
            16'd17643: data <= 8'h07;
            16'd17644: data <= 8'hE0;
            16'd17645: data <= 8'h07;
            16'd17646: data <= 8'hE0;
            16'd17647: data <= 8'h07;
            16'd17648: data <= 8'hE0;
            16'd17649: data <= 8'h07;
            16'd17650: data <= 8'hE0;
            16'd17651: data <= 8'h07;
            16'd17652: data <= 8'hE0;
            16'd17653: data <= 8'h07;
            16'd17654: data <= 8'hE0;
            16'd17655: data <= 8'h07;
            16'd17656: data <= 8'hE0;
            16'd17657: data <= 8'h07;
            16'd17658: data <= 8'hE0;
            16'd17659: data <= 8'h07;
            16'd17660: data <= 8'hE0;
            16'd17661: data <= 8'h07;
            16'd17662: data <= 8'hE0;
            16'd17663: data <= 8'h07;
            16'd17664: data <= 8'hE0;
            16'd17665: data <= 8'h07;
            16'd17666: data <= 8'hE0;
            16'd17667: data <= 8'h07;
            16'd17668: data <= 8'hE0;
            16'd17669: data <= 8'h07;
            16'd17670: data <= 8'hE0;
            16'd17671: data <= 8'h07;
            16'd17672: data <= 8'hE0;
            16'd17673: data <= 8'h07;
            16'd17674: data <= 8'hE0;
            16'd17675: data <= 8'h07;
            16'd17676: data <= 8'hE0;
            16'd17677: data <= 8'h07;
            16'd17678: data <= 8'hE0;
            16'd17679: data <= 8'h07;
            16'd17680: data <= 8'hFF;
            16'd17681: data <= 8'hFF;
            16'd17682: data <= 8'hE0;
            16'd17683: data <= 8'h07;
            16'd17684: data <= 8'hE0;
            16'd17685: data <= 8'h07;
            16'd17686: data <= 8'hE0;
            16'd17687: data <= 8'h07;
            16'd17688: data <= 8'hE0;
            16'd17689: data <= 8'h07;
            16'd17690: data <= 8'hE0;
            16'd17691: data <= 8'h07;
            16'd17692: data <= 8'hE0;
            16'd17693: data <= 8'h07;
            16'd17694: data <= 8'hE0;
            16'd17695: data <= 8'h07;
            16'd17696: data <= 8'hE0;
            16'd17697: data <= 8'h07;
            16'd17698: data <= 8'hE0;
            16'd17699: data <= 8'h07;
            16'd17700: data <= 8'hE0;
            16'd17701: data <= 8'h07;
            16'd17702: data <= 8'hE0;
            16'd17703: data <= 8'h07;
            16'd17704: data <= 8'hE0;
            16'd17705: data <= 8'h07;
            16'd17706: data <= 8'hE0;
            16'd17707: data <= 8'h07;
            16'd17708: data <= 8'hE0;
            16'd17709: data <= 8'h07;
            16'd17710: data <= 8'hE0;
            16'd17711: data <= 8'h07;
            16'd17712: data <= 8'hE0;
            16'd17713: data <= 8'h07;
            16'd17714: data <= 8'hE0;
            16'd17715: data <= 8'h07;
            16'd17716: data <= 8'hE0;
            16'd17717: data <= 8'h07;
            16'd17718: data <= 8'hE0;
            16'd17719: data <= 8'h07;
            16'd17720: data <= 8'hFF;
            16'd17721: data <= 8'hFF;
            16'd17722: data <= 8'hE0;
            16'd17723: data <= 8'h07;
            16'd17724: data <= 8'hE0;
            16'd17725: data <= 8'h07;
            16'd17726: data <= 8'hE0;
            16'd17727: data <= 8'h07;
            16'd17728: data <= 8'hE0;
            16'd17729: data <= 8'h07;
            16'd17730: data <= 8'hE0;
            16'd17731: data <= 8'h07;
            16'd17732: data <= 8'hE0;
            16'd17733: data <= 8'h07;
            16'd17734: data <= 8'hE0;
            16'd17735: data <= 8'h07;
            16'd17736: data <= 8'hE0;
            16'd17737: data <= 8'h07;
            16'd17738: data <= 8'hE0;
            16'd17739: data <= 8'h07;
            16'd17740: data <= 8'hE0;
            16'd17741: data <= 8'h07;
            16'd17742: data <= 8'hE0;
            16'd17743: data <= 8'h07;
            16'd17744: data <= 8'hE0;
            16'd17745: data <= 8'h07;
            16'd17746: data <= 8'hE0;
            16'd17747: data <= 8'h07;
            16'd17748: data <= 8'hE0;
            16'd17749: data <= 8'h07;
            16'd17750: data <= 8'hE0;
            16'd17751: data <= 8'h07;
            16'd17752: data <= 8'hE0;
            16'd17753: data <= 8'h07;
            16'd17754: data <= 8'hE0;
            16'd17755: data <= 8'h07;
            16'd17756: data <= 8'hE0;
            16'd17757: data <= 8'h07;
            16'd17758: data <= 8'hE0;
            16'd17759: data <= 8'h07;
            16'd17760: data <= 8'hFF;
            16'd17761: data <= 8'hFF;
            16'd17762: data <= 8'hE0;
            16'd17763: data <= 8'h07;
            16'd17764: data <= 8'hE0;
            16'd17765: data <= 8'h07;
            16'd17766: data <= 8'hE0;
            16'd17767: data <= 8'h07;
            16'd17768: data <= 8'hE0;
            16'd17769: data <= 8'h07;
            16'd17770: data <= 8'hE0;
            16'd17771: data <= 8'h07;
            16'd17772: data <= 8'hE0;
            16'd17773: data <= 8'h07;
            16'd17774: data <= 8'hE0;
            16'd17775: data <= 8'h07;
            16'd17776: data <= 8'hE0;
            16'd17777: data <= 8'h07;
            16'd17778: data <= 8'hE0;
            16'd17779: data <= 8'h07;
            16'd17780: data <= 8'hE0;
            16'd17781: data <= 8'h07;
            16'd17782: data <= 8'hE0;
            16'd17783: data <= 8'h07;
            16'd17784: data <= 8'hE0;
            16'd17785: data <= 8'h07;
            16'd17786: data <= 8'hE0;
            16'd17787: data <= 8'h07;
            16'd17788: data <= 8'hE0;
            16'd17789: data <= 8'h07;
            16'd17790: data <= 8'hE0;
            16'd17791: data <= 8'h07;
            16'd17792: data <= 8'hE0;
            16'd17793: data <= 8'h07;
            16'd17794: data <= 8'hE0;
            16'd17795: data <= 8'h07;
            16'd17796: data <= 8'hE0;
            16'd17797: data <= 8'h07;
            16'd17798: data <= 8'hE0;
            16'd17799: data <= 8'h07;
            16'd17800: data <= 8'hFF;
            16'd17801: data <= 8'hFF;
            16'd17802: data <= 8'hE0;
            16'd17803: data <= 8'h07;
            16'd17804: data <= 8'hE0;
            16'd17805: data <= 8'h07;
            16'd17806: data <= 8'hE0;
            16'd17807: data <= 8'h07;
            16'd17808: data <= 8'hE0;
            16'd17809: data <= 8'h07;
            16'd17810: data <= 8'hE0;
            16'd17811: data <= 8'h07;
            16'd17812: data <= 8'hE0;
            16'd17813: data <= 8'h07;
            16'd17814: data <= 8'hE0;
            16'd17815: data <= 8'h07;
            16'd17816: data <= 8'hE0;
            16'd17817: data <= 8'h07;
            16'd17818: data <= 8'hE0;
            16'd17819: data <= 8'h07;
            16'd17820: data <= 8'hE0;
            16'd17821: data <= 8'h07;
            16'd17822: data <= 8'hE0;
            16'd17823: data <= 8'h07;
            16'd17824: data <= 8'hE0;
            16'd17825: data <= 8'h07;
            16'd17826: data <= 8'hE0;
            16'd17827: data <= 8'h07;
            16'd17828: data <= 8'hE0;
            16'd17829: data <= 8'h07;
            16'd17830: data <= 8'hE0;
            16'd17831: data <= 8'h07;
            16'd17832: data <= 8'hE0;
            16'd17833: data <= 8'h07;
            16'd17834: data <= 8'hE0;
            16'd17835: data <= 8'h07;
            16'd17836: data <= 8'hE0;
            16'd17837: data <= 8'h07;
            16'd17838: data <= 8'hE0;
            16'd17839: data <= 8'h07;
            16'd17840: data <= 8'hFF;
            16'd17841: data <= 8'hFF;
            16'd17842: data <= 8'hE0;
            16'd17843: data <= 8'h07;
            16'd17844: data <= 8'hE0;
            16'd17845: data <= 8'h07;
            16'd17846: data <= 8'hE0;
            16'd17847: data <= 8'h07;
            16'd17848: data <= 8'hE0;
            16'd17849: data <= 8'h07;
            16'd17850: data <= 8'hE0;
            16'd17851: data <= 8'h07;
            16'd17852: data <= 8'hE0;
            16'd17853: data <= 8'h07;
            16'd17854: data <= 8'hE0;
            16'd17855: data <= 8'h07;
            16'd17856: data <= 8'hE0;
            16'd17857: data <= 8'h07;
            16'd17858: data <= 8'hE0;
            16'd17859: data <= 8'h07;
            16'd17860: data <= 8'hE0;
            16'd17861: data <= 8'h07;
            16'd17862: data <= 8'hE0;
            16'd17863: data <= 8'h07;
            16'd17864: data <= 8'hE0;
            16'd17865: data <= 8'h07;
            16'd17866: data <= 8'hE0;
            16'd17867: data <= 8'h07;
            16'd17868: data <= 8'hE0;
            16'd17869: data <= 8'h07;
            16'd17870: data <= 8'hE0;
            16'd17871: data <= 8'h07;
            16'd17872: data <= 8'hE0;
            16'd17873: data <= 8'h07;
            16'd17874: data <= 8'hE0;
            16'd17875: data <= 8'h07;
            16'd17876: data <= 8'hE0;
            16'd17877: data <= 8'h07;
            16'd17878: data <= 8'hE0;
            16'd17879: data <= 8'h07;
            16'd17880: data <= 8'hFF;
            16'd17881: data <= 8'hFF;
            16'd17882: data <= 8'hE0;
            16'd17883: data <= 8'h07;
            16'd17884: data <= 8'hE0;
            16'd17885: data <= 8'h07;
            16'd17886: data <= 8'hE0;
            16'd17887: data <= 8'h07;
            16'd17888: data <= 8'hE0;
            16'd17889: data <= 8'h07;
            16'd17890: data <= 8'hE0;
            16'd17891: data <= 8'h07;
            16'd17892: data <= 8'hE0;
            16'd17893: data <= 8'h07;
            16'd17894: data <= 8'hE0;
            16'd17895: data <= 8'h07;
            16'd17896: data <= 8'hE0;
            16'd17897: data <= 8'h07;
            16'd17898: data <= 8'hE0;
            16'd17899: data <= 8'h07;
            16'd17900: data <= 8'hE0;
            16'd17901: data <= 8'h07;
            16'd17902: data <= 8'hE0;
            16'd17903: data <= 8'h07;
            16'd17904: data <= 8'hE0;
            16'd17905: data <= 8'h07;
            16'd17906: data <= 8'hE0;
            16'd17907: data <= 8'h07;
            16'd17908: data <= 8'hE0;
            16'd17909: data <= 8'h07;
            16'd17910: data <= 8'hE0;
            16'd17911: data <= 8'h07;
            16'd17912: data <= 8'hE0;
            16'd17913: data <= 8'h07;
            16'd17914: data <= 8'hE0;
            16'd17915: data <= 8'h07;
            16'd17916: data <= 8'hE0;
            16'd17917: data <= 8'h07;
            16'd17918: data <= 8'hE0;
            16'd17919: data <= 8'h07;
            16'd17920: data <= 8'hFF;
            16'd17921: data <= 8'hFF;
            16'd17922: data <= 8'hE0;
            16'd17923: data <= 8'h07;
            16'd17924: data <= 8'hE0;
            16'd17925: data <= 8'h07;
            16'd17926: data <= 8'hE0;
            16'd17927: data <= 8'h07;
            16'd17928: data <= 8'hE0;
            16'd17929: data <= 8'h07;
            16'd17930: data <= 8'hE0;
            16'd17931: data <= 8'h07;
            16'd17932: data <= 8'hE0;
            16'd17933: data <= 8'h07;
            16'd17934: data <= 8'hE0;
            16'd17935: data <= 8'h07;
            16'd17936: data <= 8'hE0;
            16'd17937: data <= 8'h07;
            16'd17938: data <= 8'hE0;
            16'd17939: data <= 8'h07;
            16'd17940: data <= 8'hE0;
            16'd17941: data <= 8'h07;
            16'd17942: data <= 8'hE0;
            16'd17943: data <= 8'h07;
            16'd17944: data <= 8'hE0;
            16'd17945: data <= 8'h07;
            16'd17946: data <= 8'hE0;
            16'd17947: data <= 8'h07;
            16'd17948: data <= 8'hE0;
            16'd17949: data <= 8'h07;
            16'd17950: data <= 8'hE0;
            16'd17951: data <= 8'h07;
            16'd17952: data <= 8'hE0;
            16'd17953: data <= 8'h07;
            16'd17954: data <= 8'hE0;
            16'd17955: data <= 8'h07;
            16'd17956: data <= 8'hE0;
            16'd17957: data <= 8'h07;
            16'd17958: data <= 8'hE0;
            16'd17959: data <= 8'h07;
            16'd17960: data <= 8'hFF;
            16'd17961: data <= 8'hFF;
            16'd17962: data <= 8'hE0;
            16'd17963: data <= 8'h07;
            16'd17964: data <= 8'hE0;
            16'd17965: data <= 8'h07;
            16'd17966: data <= 8'hE0;
            16'd17967: data <= 8'h07;
            16'd17968: data <= 8'hE0;
            16'd17969: data <= 8'h07;
            16'd17970: data <= 8'hE0;
            16'd17971: data <= 8'h07;
            16'd17972: data <= 8'hE0;
            16'd17973: data <= 8'h07;
            16'd17974: data <= 8'hE0;
            16'd17975: data <= 8'h07;
            16'd17976: data <= 8'hE0;
            16'd17977: data <= 8'h07;
            16'd17978: data <= 8'hE0;
            16'd17979: data <= 8'h07;
            16'd17980: data <= 8'hE0;
            16'd17981: data <= 8'h07;
            16'd17982: data <= 8'hE0;
            16'd17983: data <= 8'h07;
            16'd17984: data <= 8'hE0;
            16'd17985: data <= 8'h07;
            16'd17986: data <= 8'hE0;
            16'd17987: data <= 8'h07;
            16'd17988: data <= 8'hE0;
            16'd17989: data <= 8'h07;
            16'd17990: data <= 8'hE0;
            16'd17991: data <= 8'h07;
            16'd17992: data <= 8'hE0;
            16'd17993: data <= 8'h07;
            16'd17994: data <= 8'hE0;
            16'd17995: data <= 8'h07;
            16'd17996: data <= 8'hE0;
            16'd17997: data <= 8'h07;
            16'd17998: data <= 8'hE0;
            16'd17999: data <= 8'h07;
            16'd18000: data <= 8'hFF;
            16'd18001: data <= 8'hFF;
            16'd18002: data <= 8'hE0;
            16'd18003: data <= 8'h07;
            16'd18004: data <= 8'hE0;
            16'd18005: data <= 8'h07;
            16'd18006: data <= 8'hE0;
            16'd18007: data <= 8'h07;
            16'd18008: data <= 8'hE0;
            16'd18009: data <= 8'h07;
            16'd18010: data <= 8'hE0;
            16'd18011: data <= 8'h07;
            16'd18012: data <= 8'hE0;
            16'd18013: data <= 8'h07;
            16'd18014: data <= 8'hE0;
            16'd18015: data <= 8'h07;
            16'd18016: data <= 8'hE0;
            16'd18017: data <= 8'h07;
            16'd18018: data <= 8'hE0;
            16'd18019: data <= 8'h07;
            16'd18020: data <= 8'hE0;
            16'd18021: data <= 8'h07;
            16'd18022: data <= 8'hE0;
            16'd18023: data <= 8'h07;
            16'd18024: data <= 8'hE0;
            16'd18025: data <= 8'h07;
            16'd18026: data <= 8'hE0;
            16'd18027: data <= 8'h07;
            16'd18028: data <= 8'hE0;
            16'd18029: data <= 8'h07;
            16'd18030: data <= 8'hE0;
            16'd18031: data <= 8'h07;
            16'd18032: data <= 8'hE0;
            16'd18033: data <= 8'h07;
            16'd18034: data <= 8'hE0;
            16'd18035: data <= 8'h07;
            16'd18036: data <= 8'hE0;
            16'd18037: data <= 8'h07;
            16'd18038: data <= 8'hE0;
            16'd18039: data <= 8'h07;
            16'd18040: data <= 8'hFF;
            16'd18041: data <= 8'hFF;
            16'd18042: data <= 8'hE0;
            16'd18043: data <= 8'h07;
            16'd18044: data <= 8'hE0;
            16'd18045: data <= 8'h07;
            16'd18046: data <= 8'hE0;
            16'd18047: data <= 8'h07;
            16'd18048: data <= 8'hE0;
            16'd18049: data <= 8'h07;
            16'd18050: data <= 8'hE0;
            16'd18051: data <= 8'h07;
            16'd18052: data <= 8'hE0;
            16'd18053: data <= 8'h07;
            16'd18054: data <= 8'hE0;
            16'd18055: data <= 8'h07;
            16'd18056: data <= 8'hE0;
            16'd18057: data <= 8'h07;
            16'd18058: data <= 8'hE0;
            16'd18059: data <= 8'h07;
            16'd18060: data <= 8'hE0;
            16'd18061: data <= 8'h07;
            16'd18062: data <= 8'hE0;
            16'd18063: data <= 8'h07;
            16'd18064: data <= 8'hE0;
            16'd18065: data <= 8'h07;
            16'd18066: data <= 8'hE0;
            16'd18067: data <= 8'h07;
            16'd18068: data <= 8'hE0;
            16'd18069: data <= 8'h07;
            16'd18070: data <= 8'hE0;
            16'd18071: data <= 8'h07;
            16'd18072: data <= 8'hE0;
            16'd18073: data <= 8'h07;
            16'd18074: data <= 8'hE0;
            16'd18075: data <= 8'h07;
            16'd18076: data <= 8'hE0;
            16'd18077: data <= 8'h07;
            16'd18078: data <= 8'hE0;
            16'd18079: data <= 8'h07;
            16'd18080: data <= 8'hFF;
            16'd18081: data <= 8'hFF;
            16'd18082: data <= 8'hE0;
            16'd18083: data <= 8'h07;
            16'd18084: data <= 8'hE0;
            16'd18085: data <= 8'h07;
            16'd18086: data <= 8'hE0;
            16'd18087: data <= 8'h07;
            16'd18088: data <= 8'hE0;
            16'd18089: data <= 8'h07;
            16'd18090: data <= 8'hE0;
            16'd18091: data <= 8'h07;
            16'd18092: data <= 8'hE0;
            16'd18093: data <= 8'h07;
            16'd18094: data <= 8'hE0;
            16'd18095: data <= 8'h07;
            16'd18096: data <= 8'hE0;
            16'd18097: data <= 8'h07;
            16'd18098: data <= 8'hE0;
            16'd18099: data <= 8'h07;
            16'd18100: data <= 8'hE0;
            16'd18101: data <= 8'h07;
            16'd18102: data <= 8'hE0;
            16'd18103: data <= 8'h07;
            16'd18104: data <= 8'hE0;
            16'd18105: data <= 8'h07;
            16'd18106: data <= 8'hE0;
            16'd18107: data <= 8'h07;
            16'd18108: data <= 8'hE0;
            16'd18109: data <= 8'h07;
            16'd18110: data <= 8'hE0;
            16'd18111: data <= 8'h07;
            16'd18112: data <= 8'hE0;
            16'd18113: data <= 8'h07;
            16'd18114: data <= 8'hE0;
            16'd18115: data <= 8'h07;
            16'd18116: data <= 8'hE0;
            16'd18117: data <= 8'h07;
            16'd18118: data <= 8'hE0;
            16'd18119: data <= 8'h07;
            16'd18120: data <= 8'hFF;
            16'd18121: data <= 8'hFF;
            16'd18122: data <= 8'hE0;
            16'd18123: data <= 8'h07;
            16'd18124: data <= 8'hE0;
            16'd18125: data <= 8'h07;
            16'd18126: data <= 8'hE0;
            16'd18127: data <= 8'h07;
            16'd18128: data <= 8'hE0;
            16'd18129: data <= 8'h07;
            16'd18130: data <= 8'hE0;
            16'd18131: data <= 8'h07;
            16'd18132: data <= 8'hE0;
            16'd18133: data <= 8'h07;
            16'd18134: data <= 8'hE0;
            16'd18135: data <= 8'h07;
            16'd18136: data <= 8'hE0;
            16'd18137: data <= 8'h07;
            16'd18138: data <= 8'hE0;
            16'd18139: data <= 8'h07;
            16'd18140: data <= 8'hE0;
            16'd18141: data <= 8'h07;
            16'd18142: data <= 8'hE0;
            16'd18143: data <= 8'h07;
            16'd18144: data <= 8'hE0;
            16'd18145: data <= 8'h07;
            16'd18146: data <= 8'hE0;
            16'd18147: data <= 8'h07;
            16'd18148: data <= 8'hE0;
            16'd18149: data <= 8'h07;
            16'd18150: data <= 8'hE0;
            16'd18151: data <= 8'h07;
            16'd18152: data <= 8'hE0;
            16'd18153: data <= 8'h07;
            16'd18154: data <= 8'hE0;
            16'd18155: data <= 8'h07;
            16'd18156: data <= 8'hE0;
            16'd18157: data <= 8'h07;
            16'd18158: data <= 8'hE0;
            16'd18159: data <= 8'h07;
            16'd18160: data <= 8'hFF;
            16'd18161: data <= 8'hFF;
            16'd18162: data <= 8'hE0;
            16'd18163: data <= 8'h07;
            16'd18164: data <= 8'hE0;
            16'd18165: data <= 8'h07;
            16'd18166: data <= 8'hE0;
            16'd18167: data <= 8'h07;
            16'd18168: data <= 8'hE0;
            16'd18169: data <= 8'h07;
            16'd18170: data <= 8'hE0;
            16'd18171: data <= 8'h07;
            16'd18172: data <= 8'hE0;
            16'd18173: data <= 8'h07;
            16'd18174: data <= 8'hE0;
            16'd18175: data <= 8'h07;
            16'd18176: data <= 8'hE0;
            16'd18177: data <= 8'h07;
            16'd18178: data <= 8'hE0;
            16'd18179: data <= 8'h07;
            16'd18180: data <= 8'hE0;
            16'd18181: data <= 8'h07;
            16'd18182: data <= 8'hE0;
            16'd18183: data <= 8'h07;
            16'd18184: data <= 8'hE0;
            16'd18185: data <= 8'h07;
            16'd18186: data <= 8'hE0;
            16'd18187: data <= 8'h07;
            16'd18188: data <= 8'hE0;
            16'd18189: data <= 8'h07;
            16'd18190: data <= 8'hE0;
            16'd18191: data <= 8'h07;
            16'd18192: data <= 8'hE0;
            16'd18193: data <= 8'h07;
            16'd18194: data <= 8'hE0;
            16'd18195: data <= 8'h07;
            16'd18196: data <= 8'hE0;
            16'd18197: data <= 8'h07;
            16'd18198: data <= 8'hE0;
            16'd18199: data <= 8'h07;
            16'd18200: data <= 8'hFF;
            16'd18201: data <= 8'hFF;
            16'd18202: data <= 8'hE0;
            16'd18203: data <= 8'h07;
            16'd18204: data <= 8'hE0;
            16'd18205: data <= 8'h07;
            16'd18206: data <= 8'hE0;
            16'd18207: data <= 8'h07;
            16'd18208: data <= 8'hE0;
            16'd18209: data <= 8'h07;
            16'd18210: data <= 8'hE0;
            16'd18211: data <= 8'h07;
            16'd18212: data <= 8'hE0;
            16'd18213: data <= 8'h07;
            16'd18214: data <= 8'hE0;
            16'd18215: data <= 8'h07;
            16'd18216: data <= 8'hE0;
            16'd18217: data <= 8'h07;
            16'd18218: data <= 8'hE0;
            16'd18219: data <= 8'h07;
            16'd18220: data <= 8'hE0;
            16'd18221: data <= 8'h07;
            16'd18222: data <= 8'hE0;
            16'd18223: data <= 8'h07;
            16'd18224: data <= 8'hE0;
            16'd18225: data <= 8'h07;
            16'd18226: data <= 8'hE0;
            16'd18227: data <= 8'h07;
            16'd18228: data <= 8'hE0;
            16'd18229: data <= 8'h07;
            16'd18230: data <= 8'hE0;
            16'd18231: data <= 8'h07;
            16'd18232: data <= 8'hE0;
            16'd18233: data <= 8'h07;
            16'd18234: data <= 8'hE0;
            16'd18235: data <= 8'h07;
            16'd18236: data <= 8'hE0;
            16'd18237: data <= 8'h07;
            16'd18238: data <= 8'hE0;
            16'd18239: data <= 8'h07;
            16'd18240: data <= 8'hFF;
            16'd18241: data <= 8'hFF;
            16'd18242: data <= 8'hE0;
            16'd18243: data <= 8'h07;
            16'd18244: data <= 8'hE0;
            16'd18245: data <= 8'h07;
            16'd18246: data <= 8'hE0;
            16'd18247: data <= 8'h07;
            16'd18248: data <= 8'hE0;
            16'd18249: data <= 8'h07;
            16'd18250: data <= 8'hE0;
            16'd18251: data <= 8'h07;
            16'd18252: data <= 8'hE0;
            16'd18253: data <= 8'h07;
            16'd18254: data <= 8'hE0;
            16'd18255: data <= 8'h07;
            16'd18256: data <= 8'hE0;
            16'd18257: data <= 8'h07;
            16'd18258: data <= 8'hE0;
            16'd18259: data <= 8'h07;
            16'd18260: data <= 8'hE0;
            16'd18261: data <= 8'h07;
            16'd18262: data <= 8'hE0;
            16'd18263: data <= 8'h07;
            16'd18264: data <= 8'hE0;
            16'd18265: data <= 8'h07;
            16'd18266: data <= 8'hE0;
            16'd18267: data <= 8'h07;
            16'd18268: data <= 8'hE0;
            16'd18269: data <= 8'h07;
            16'd18270: data <= 8'hE0;
            16'd18271: data <= 8'h07;
            16'd18272: data <= 8'hE0;
            16'd18273: data <= 8'h07;
            16'd18274: data <= 8'hE0;
            16'd18275: data <= 8'h07;
            16'd18276: data <= 8'hE0;
            16'd18277: data <= 8'h07;
            16'd18278: data <= 8'hE0;
            16'd18279: data <= 8'h07;
            16'd18280: data <= 8'hFF;
            16'd18281: data <= 8'hFF;
            16'd18282: data <= 8'hE0;
            16'd18283: data <= 8'h07;
            16'd18284: data <= 8'hE0;
            16'd18285: data <= 8'h07;
            16'd18286: data <= 8'hE0;
            16'd18287: data <= 8'h07;
            16'd18288: data <= 8'hE0;
            16'd18289: data <= 8'h07;
            16'd18290: data <= 8'hE0;
            16'd18291: data <= 8'h07;
            16'd18292: data <= 8'hE0;
            16'd18293: data <= 8'h07;
            16'd18294: data <= 8'hE0;
            16'd18295: data <= 8'h07;
            16'd18296: data <= 8'hE0;
            16'd18297: data <= 8'h07;
            16'd18298: data <= 8'hE0;
            16'd18299: data <= 8'h07;
            16'd18300: data <= 8'hE0;
            16'd18301: data <= 8'h07;
            16'd18302: data <= 8'hE0;
            16'd18303: data <= 8'h07;
            16'd18304: data <= 8'hE0;
            16'd18305: data <= 8'h07;
            16'd18306: data <= 8'hE0;
            16'd18307: data <= 8'h07;
            16'd18308: data <= 8'hE0;
            16'd18309: data <= 8'h07;
            16'd18310: data <= 8'hE0;
            16'd18311: data <= 8'h07;
            16'd18312: data <= 8'hE0;
            16'd18313: data <= 8'h07;
            16'd18314: data <= 8'hE0;
            16'd18315: data <= 8'h07;
            16'd18316: data <= 8'hE0;
            16'd18317: data <= 8'h07;
            16'd18318: data <= 8'hE0;
            16'd18319: data <= 8'h07;
            16'd18320: data <= 8'hFF;
            16'd18321: data <= 8'hFF;
            16'd18322: data <= 8'hE0;
            16'd18323: data <= 8'h07;
            16'd18324: data <= 8'hE0;
            16'd18325: data <= 8'h07;
            16'd18326: data <= 8'hE0;
            16'd18327: data <= 8'h07;
            16'd18328: data <= 8'hE0;
            16'd18329: data <= 8'h07;
            16'd18330: data <= 8'hE0;
            16'd18331: data <= 8'h07;
            16'd18332: data <= 8'hE0;
            16'd18333: data <= 8'h07;
            16'd18334: data <= 8'hE0;
            16'd18335: data <= 8'h07;
            16'd18336: data <= 8'hE0;
            16'd18337: data <= 8'h07;
            16'd18338: data <= 8'hE0;
            16'd18339: data <= 8'h07;
            16'd18340: data <= 8'hE0;
            16'd18341: data <= 8'h07;
            16'd18342: data <= 8'hE0;
            16'd18343: data <= 8'h07;
            16'd18344: data <= 8'hE0;
            16'd18345: data <= 8'h07;
            16'd18346: data <= 8'hE0;
            16'd18347: data <= 8'h07;
            16'd18348: data <= 8'hE0;
            16'd18349: data <= 8'h07;
            16'd18350: data <= 8'hE0;
            16'd18351: data <= 8'h07;
            16'd18352: data <= 8'hE0;
            16'd18353: data <= 8'h07;
            16'd18354: data <= 8'hE0;
            16'd18355: data <= 8'h07;
            16'd18356: data <= 8'hE0;
            16'd18357: data <= 8'h07;
            16'd18358: data <= 8'hE0;
            16'd18359: data <= 8'h07;
            16'd18360: data <= 8'hFF;
            16'd18361: data <= 8'hFF;
            16'd18362: data <= 8'hE0;
            16'd18363: data <= 8'h07;
            16'd18364: data <= 8'hE0;
            16'd18365: data <= 8'h07;
            16'd18366: data <= 8'hE0;
            16'd18367: data <= 8'h07;
            16'd18368: data <= 8'hE0;
            16'd18369: data <= 8'h07;
            16'd18370: data <= 8'hE0;
            16'd18371: data <= 8'h07;
            16'd18372: data <= 8'hE0;
            16'd18373: data <= 8'h07;
            16'd18374: data <= 8'hE0;
            16'd18375: data <= 8'h07;
            16'd18376: data <= 8'hE0;
            16'd18377: data <= 8'h07;
            16'd18378: data <= 8'hE0;
            16'd18379: data <= 8'h07;
            16'd18380: data <= 8'hE0;
            16'd18381: data <= 8'h07;
            16'd18382: data <= 8'hE0;
            16'd18383: data <= 8'h07;
            16'd18384: data <= 8'hE0;
            16'd18385: data <= 8'h07;
            16'd18386: data <= 8'hE0;
            16'd18387: data <= 8'h07;
            16'd18388: data <= 8'hE0;
            16'd18389: data <= 8'h07;
            16'd18390: data <= 8'hE0;
            16'd18391: data <= 8'h07;
            16'd18392: data <= 8'hE0;
            16'd18393: data <= 8'h07;
            16'd18394: data <= 8'hE0;
            16'd18395: data <= 8'h07;
            16'd18396: data <= 8'hE0;
            16'd18397: data <= 8'h07;
            16'd18398: data <= 8'hE0;
            16'd18399: data <= 8'h07;
            16'd18400: data <= 8'hFF;
            16'd18401: data <= 8'hFF;
            16'd18402: data <= 8'hE0;
            16'd18403: data <= 8'h07;
            16'd18404: data <= 8'hE0;
            16'd18405: data <= 8'h07;
            16'd18406: data <= 8'hE0;
            16'd18407: data <= 8'h07;
            16'd18408: data <= 8'hE0;
            16'd18409: data <= 8'h07;
            16'd18410: data <= 8'hE0;
            16'd18411: data <= 8'h07;
            16'd18412: data <= 8'hE0;
            16'd18413: data <= 8'h07;
            16'd18414: data <= 8'hE0;
            16'd18415: data <= 8'h07;
            16'd18416: data <= 8'hE0;
            16'd18417: data <= 8'h07;
            16'd18418: data <= 8'hE0;
            16'd18419: data <= 8'h07;
            16'd18420: data <= 8'hE0;
            16'd18421: data <= 8'h07;
            16'd18422: data <= 8'hE0;
            16'd18423: data <= 8'h07;
            16'd18424: data <= 8'hE0;
            16'd18425: data <= 8'h07;
            16'd18426: data <= 8'hE0;
            16'd18427: data <= 8'h07;
            16'd18428: data <= 8'hE0;
            16'd18429: data <= 8'h07;
            16'd18430: data <= 8'hE0;
            16'd18431: data <= 8'h07;
            16'd18432: data <= 8'hE0;
            16'd18433: data <= 8'h07;
            16'd18434: data <= 8'hE0;
            16'd18435: data <= 8'h07;
            16'd18436: data <= 8'hE0;
            16'd18437: data <= 8'h07;
            16'd18438: data <= 8'hE0;
            16'd18439: data <= 8'h07;
            16'd18440: data <= 8'hFF;
            16'd18441: data <= 8'hFF;
            16'd18442: data <= 8'hE0;
            16'd18443: data <= 8'h07;
            16'd18444: data <= 8'hE0;
            16'd18445: data <= 8'h07;
            16'd18446: data <= 8'hE0;
            16'd18447: data <= 8'h07;
            16'd18448: data <= 8'hE0;
            16'd18449: data <= 8'h07;
            16'd18450: data <= 8'hE0;
            16'd18451: data <= 8'h07;
            16'd18452: data <= 8'hE0;
            16'd18453: data <= 8'h07;
            16'd18454: data <= 8'hE0;
            16'd18455: data <= 8'h07;
            16'd18456: data <= 8'hE0;
            16'd18457: data <= 8'h07;
            16'd18458: data <= 8'hE0;
            16'd18459: data <= 8'h07;
            16'd18460: data <= 8'hE0;
            16'd18461: data <= 8'h07;
            16'd18462: data <= 8'hE0;
            16'd18463: data <= 8'h07;
            16'd18464: data <= 8'hE0;
            16'd18465: data <= 8'h07;
            16'd18466: data <= 8'hE0;
            16'd18467: data <= 8'h07;
            16'd18468: data <= 8'hE0;
            16'd18469: data <= 8'h07;
            16'd18470: data <= 8'hE0;
            16'd18471: data <= 8'h07;
            16'd18472: data <= 8'hE0;
            16'd18473: data <= 8'h07;
            16'd18474: data <= 8'hE0;
            16'd18475: data <= 8'h07;
            16'd18476: data <= 8'hE0;
            16'd18477: data <= 8'h07;
            16'd18478: data <= 8'hE0;
            16'd18479: data <= 8'h07;
            16'd18480: data <= 8'hFF;
            16'd18481: data <= 8'hFF;
            16'd18482: data <= 8'hE0;
            16'd18483: data <= 8'h07;
            16'd18484: data <= 8'hE0;
            16'd18485: data <= 8'h07;
            16'd18486: data <= 8'hE0;
            16'd18487: data <= 8'h07;
            16'd18488: data <= 8'hE0;
            16'd18489: data <= 8'h07;
            16'd18490: data <= 8'hE0;
            16'd18491: data <= 8'h07;
            16'd18492: data <= 8'hE0;
            16'd18493: data <= 8'h07;
            16'd18494: data <= 8'hE0;
            16'd18495: data <= 8'h07;
            16'd18496: data <= 8'hE0;
            16'd18497: data <= 8'h07;
            16'd18498: data <= 8'hE0;
            16'd18499: data <= 8'h07;
            16'd18500: data <= 8'hE0;
            16'd18501: data <= 8'h07;
            16'd18502: data <= 8'hE0;
            16'd18503: data <= 8'h07;
            16'd18504: data <= 8'hE0;
            16'd18505: data <= 8'h07;
            16'd18506: data <= 8'hE0;
            16'd18507: data <= 8'h07;
            16'd18508: data <= 8'hE0;
            16'd18509: data <= 8'h07;
            16'd18510: data <= 8'hE0;
            16'd18511: data <= 8'h07;
            16'd18512: data <= 8'hE0;
            16'd18513: data <= 8'h07;
            16'd18514: data <= 8'hE0;
            16'd18515: data <= 8'h07;
            16'd18516: data <= 8'hE0;
            16'd18517: data <= 8'h07;
            16'd18518: data <= 8'hE0;
            16'd18519: data <= 8'h07;
            16'd18520: data <= 8'hFF;
            16'd18521: data <= 8'hFF;
            16'd18522: data <= 8'hE0;
            16'd18523: data <= 8'h07;
            16'd18524: data <= 8'hE0;
            16'd18525: data <= 8'h07;
            16'd18526: data <= 8'hE0;
            16'd18527: data <= 8'h07;
            16'd18528: data <= 8'hE0;
            16'd18529: data <= 8'h07;
            16'd18530: data <= 8'hE0;
            16'd18531: data <= 8'h07;
            16'd18532: data <= 8'hE0;
            16'd18533: data <= 8'h07;
            16'd18534: data <= 8'hE0;
            16'd18535: data <= 8'h07;
            16'd18536: data <= 8'hE0;
            16'd18537: data <= 8'h07;
            16'd18538: data <= 8'hE0;
            16'd18539: data <= 8'h07;
            16'd18540: data <= 8'hE0;
            16'd18541: data <= 8'h07;
            16'd18542: data <= 8'hE0;
            16'd18543: data <= 8'h07;
            16'd18544: data <= 8'hE0;
            16'd18545: data <= 8'h07;
            16'd18546: data <= 8'hE0;
            16'd18547: data <= 8'h07;
            16'd18548: data <= 8'hE0;
            16'd18549: data <= 8'h07;
            16'd18550: data <= 8'hE0;
            16'd18551: data <= 8'h07;
            16'd18552: data <= 8'hE0;
            16'd18553: data <= 8'h07;
            16'd18554: data <= 8'hE0;
            16'd18555: data <= 8'h07;
            16'd18556: data <= 8'hE0;
            16'd18557: data <= 8'h07;
            16'd18558: data <= 8'hE0;
            16'd18559: data <= 8'h07;
            16'd18560: data <= 8'hFF;
            16'd18561: data <= 8'hFF;
            16'd18562: data <= 8'hE0;
            16'd18563: data <= 8'h07;
            16'd18564: data <= 8'hE0;
            16'd18565: data <= 8'h07;
            16'd18566: data <= 8'hE0;
            16'd18567: data <= 8'h07;
            16'd18568: data <= 8'hE0;
            16'd18569: data <= 8'h07;
            16'd18570: data <= 8'hE0;
            16'd18571: data <= 8'h07;
            16'd18572: data <= 8'hE0;
            16'd18573: data <= 8'h07;
            16'd18574: data <= 8'hE0;
            16'd18575: data <= 8'h07;
            16'd18576: data <= 8'hE0;
            16'd18577: data <= 8'h07;
            16'd18578: data <= 8'hE0;
            16'd18579: data <= 8'h07;
            16'd18580: data <= 8'hE0;
            16'd18581: data <= 8'h07;
            16'd18582: data <= 8'hE0;
            16'd18583: data <= 8'h07;
            16'd18584: data <= 8'hE0;
            16'd18585: data <= 8'h07;
            16'd18586: data <= 8'hE0;
            16'd18587: data <= 8'h07;
            16'd18588: data <= 8'hE0;
            16'd18589: data <= 8'h07;
            16'd18590: data <= 8'hE0;
            16'd18591: data <= 8'h07;
            16'd18592: data <= 8'hE0;
            16'd18593: data <= 8'h07;
            16'd18594: data <= 8'hE0;
            16'd18595: data <= 8'h07;
            16'd18596: data <= 8'hE0;
            16'd18597: data <= 8'h07;
            16'd18598: data <= 8'hE0;
            16'd18599: data <= 8'h07;
            16'd18600: data <= 8'hFF;
            16'd18601: data <= 8'hFF;
            16'd18602: data <= 8'hE0;
            16'd18603: data <= 8'h07;
            16'd18604: data <= 8'hE0;
            16'd18605: data <= 8'h07;
            16'd18606: data <= 8'hE0;
            16'd18607: data <= 8'h07;
            16'd18608: data <= 8'hE0;
            16'd18609: data <= 8'h07;
            16'd18610: data <= 8'hE0;
            16'd18611: data <= 8'h07;
            16'd18612: data <= 8'hE0;
            16'd18613: data <= 8'h07;
            16'd18614: data <= 8'hE0;
            16'd18615: data <= 8'h07;
            16'd18616: data <= 8'hE0;
            16'd18617: data <= 8'h07;
            16'd18618: data <= 8'hE0;
            16'd18619: data <= 8'h07;
            16'd18620: data <= 8'hE0;
            16'd18621: data <= 8'h07;
            16'd18622: data <= 8'hE0;
            16'd18623: data <= 8'h07;
            16'd18624: data <= 8'hE0;
            16'd18625: data <= 8'h07;
            16'd18626: data <= 8'hE0;
            16'd18627: data <= 8'h07;
            16'd18628: data <= 8'hE0;
            16'd18629: data <= 8'h07;
            16'd18630: data <= 8'hE0;
            16'd18631: data <= 8'h07;
            16'd18632: data <= 8'hE0;
            16'd18633: data <= 8'h07;
            16'd18634: data <= 8'hE0;
            16'd18635: data <= 8'h07;
            16'd18636: data <= 8'hE0;
            16'd18637: data <= 8'h07;
            16'd18638: data <= 8'hE0;
            16'd18639: data <= 8'h07;
            16'd18640: data <= 8'hFF;
            16'd18641: data <= 8'hFF;
            16'd18642: data <= 8'hE0;
            16'd18643: data <= 8'h07;
            16'd18644: data <= 8'hE0;
            16'd18645: data <= 8'h07;
            16'd18646: data <= 8'hE0;
            16'd18647: data <= 8'h07;
            16'd18648: data <= 8'hE0;
            16'd18649: data <= 8'h07;
            16'd18650: data <= 8'hE0;
            16'd18651: data <= 8'h07;
            16'd18652: data <= 8'hE0;
            16'd18653: data <= 8'h07;
            16'd18654: data <= 8'hE0;
            16'd18655: data <= 8'h07;
            16'd18656: data <= 8'hE0;
            16'd18657: data <= 8'h07;
            16'd18658: data <= 8'hE0;
            16'd18659: data <= 8'h07;
            16'd18660: data <= 8'hE0;
            16'd18661: data <= 8'h07;
            16'd18662: data <= 8'hE0;
            16'd18663: data <= 8'h07;
            16'd18664: data <= 8'hE0;
            16'd18665: data <= 8'h07;
            16'd18666: data <= 8'hE0;
            16'd18667: data <= 8'h07;
            16'd18668: data <= 8'hE0;
            16'd18669: data <= 8'h07;
            16'd18670: data <= 8'hE0;
            16'd18671: data <= 8'h07;
            16'd18672: data <= 8'hE0;
            16'd18673: data <= 8'h07;
            16'd18674: data <= 8'hE0;
            16'd18675: data <= 8'h07;
            16'd18676: data <= 8'hE0;
            16'd18677: data <= 8'h07;
            16'd18678: data <= 8'hE0;
            16'd18679: data <= 8'h07;
            16'd18680: data <= 8'hFF;
            16'd18681: data <= 8'hFF;
            16'd18682: data <= 8'hE0;
            16'd18683: data <= 8'h07;
            16'd18684: data <= 8'hE0;
            16'd18685: data <= 8'h07;
            16'd18686: data <= 8'hE0;
            16'd18687: data <= 8'h07;
            16'd18688: data <= 8'hE0;
            16'd18689: data <= 8'h07;
            16'd18690: data <= 8'hE0;
            16'd18691: data <= 8'h07;
            16'd18692: data <= 8'hE0;
            16'd18693: data <= 8'h07;
            16'd18694: data <= 8'hE0;
            16'd18695: data <= 8'h07;
            16'd18696: data <= 8'hE0;
            16'd18697: data <= 8'h07;
            16'd18698: data <= 8'hE0;
            16'd18699: data <= 8'h07;
            16'd18700: data <= 8'hE0;
            16'd18701: data <= 8'h07;
            16'd18702: data <= 8'hE0;
            16'd18703: data <= 8'h07;
            16'd18704: data <= 8'hE0;
            16'd18705: data <= 8'h07;
            16'd18706: data <= 8'hE0;
            16'd18707: data <= 8'h07;
            16'd18708: data <= 8'hE0;
            16'd18709: data <= 8'h07;
            16'd18710: data <= 8'hE0;
            16'd18711: data <= 8'h07;
            16'd18712: data <= 8'hE0;
            16'd18713: data <= 8'h07;
            16'd18714: data <= 8'hE0;
            16'd18715: data <= 8'h07;
            16'd18716: data <= 8'hE0;
            16'd18717: data <= 8'h07;
            16'd18718: data <= 8'hE0;
            16'd18719: data <= 8'h07;
            16'd18720: data <= 8'hFF;
            16'd18721: data <= 8'hFF;
            16'd18722: data <= 8'hE0;
            16'd18723: data <= 8'h07;
            16'd18724: data <= 8'hE0;
            16'd18725: data <= 8'h07;
            16'd18726: data <= 8'hE0;
            16'd18727: data <= 8'h07;
            16'd18728: data <= 8'hE0;
            16'd18729: data <= 8'h07;
            16'd18730: data <= 8'hE0;
            16'd18731: data <= 8'h07;
            16'd18732: data <= 8'hE0;
            16'd18733: data <= 8'h07;
            16'd18734: data <= 8'hE0;
            16'd18735: data <= 8'h07;
            16'd18736: data <= 8'hE0;
            16'd18737: data <= 8'h07;
            16'd18738: data <= 8'hE0;
            16'd18739: data <= 8'h07;
            16'd18740: data <= 8'hE0;
            16'd18741: data <= 8'h07;
            16'd18742: data <= 8'hE0;
            16'd18743: data <= 8'h07;
            16'd18744: data <= 8'hE0;
            16'd18745: data <= 8'h07;
            16'd18746: data <= 8'hE0;
            16'd18747: data <= 8'h07;
            16'd18748: data <= 8'hE0;
            16'd18749: data <= 8'h07;
            16'd18750: data <= 8'hE0;
            16'd18751: data <= 8'h07;
            16'd18752: data <= 8'hE0;
            16'd18753: data <= 8'h07;
            16'd18754: data <= 8'hE0;
            16'd18755: data <= 8'h07;
            16'd18756: data <= 8'hE0;
            16'd18757: data <= 8'h07;
            16'd18758: data <= 8'hE0;
            16'd18759: data <= 8'h07;
            16'd18760: data <= 8'hFF;
            16'd18761: data <= 8'hFF;
            16'd18762: data <= 8'hE0;
            16'd18763: data <= 8'h07;
            16'd18764: data <= 8'hE0;
            16'd18765: data <= 8'h07;
            16'd18766: data <= 8'hE0;
            16'd18767: data <= 8'h07;
            16'd18768: data <= 8'hE0;
            16'd18769: data <= 8'h07;
            16'd18770: data <= 8'hE0;
            16'd18771: data <= 8'h07;
            16'd18772: data <= 8'hE0;
            16'd18773: data <= 8'h07;
            16'd18774: data <= 8'hE0;
            16'd18775: data <= 8'h07;
            16'd18776: data <= 8'hE0;
            16'd18777: data <= 8'h07;
            16'd18778: data <= 8'hE0;
            16'd18779: data <= 8'h07;
            16'd18780: data <= 8'hE0;
            16'd18781: data <= 8'h07;
            16'd18782: data <= 8'hE0;
            16'd18783: data <= 8'h07;
            16'd18784: data <= 8'hE0;
            16'd18785: data <= 8'h07;
            16'd18786: data <= 8'hE0;
            16'd18787: data <= 8'h07;
            16'd18788: data <= 8'hE0;
            16'd18789: data <= 8'h07;
            16'd18790: data <= 8'hE0;
            16'd18791: data <= 8'h07;
            16'd18792: data <= 8'hE0;
            16'd18793: data <= 8'h07;
            16'd18794: data <= 8'hE0;
            16'd18795: data <= 8'h07;
            16'd18796: data <= 8'hE0;
            16'd18797: data <= 8'h07;
            16'd18798: data <= 8'hE0;
            16'd18799: data <= 8'h07;
            16'd18800: data <= 8'hFF;
            16'd18801: data <= 8'hFF;
            16'd18802: data <= 8'hE0;
            16'd18803: data <= 8'h07;
            16'd18804: data <= 8'hE0;
            16'd18805: data <= 8'h07;
            16'd18806: data <= 8'hE0;
            16'd18807: data <= 8'h07;
            16'd18808: data <= 8'hE0;
            16'd18809: data <= 8'h07;
            16'd18810: data <= 8'hE0;
            16'd18811: data <= 8'h07;
            16'd18812: data <= 8'hE0;
            16'd18813: data <= 8'h07;
            16'd18814: data <= 8'hE0;
            16'd18815: data <= 8'h07;
            16'd18816: data <= 8'hE0;
            16'd18817: data <= 8'h07;
            16'd18818: data <= 8'hE0;
            16'd18819: data <= 8'h07;
            16'd18820: data <= 8'hE0;
            16'd18821: data <= 8'h07;
            16'd18822: data <= 8'hE0;
            16'd18823: data <= 8'h07;
            16'd18824: data <= 8'hE0;
            16'd18825: data <= 8'h07;
            16'd18826: data <= 8'hE0;
            16'd18827: data <= 8'h07;
            16'd18828: data <= 8'hE0;
            16'd18829: data <= 8'h07;
            16'd18830: data <= 8'hE0;
            16'd18831: data <= 8'h07;
            16'd18832: data <= 8'hE0;
            16'd18833: data <= 8'h07;
            16'd18834: data <= 8'hE0;
            16'd18835: data <= 8'h07;
            16'd18836: data <= 8'hE0;
            16'd18837: data <= 8'h07;
            16'd18838: data <= 8'hE0;
            16'd18839: data <= 8'h07;
            16'd18840: data <= 8'hFF;
            16'd18841: data <= 8'hFF;
            16'd18842: data <= 8'hE0;
            16'd18843: data <= 8'h07;
            16'd18844: data <= 8'hE0;
            16'd18845: data <= 8'h07;
            16'd18846: data <= 8'hE0;
            16'd18847: data <= 8'h07;
            16'd18848: data <= 8'hE0;
            16'd18849: data <= 8'h07;
            16'd18850: data <= 8'hE0;
            16'd18851: data <= 8'h07;
            16'd18852: data <= 8'hE0;
            16'd18853: data <= 8'h07;
            16'd18854: data <= 8'hE0;
            16'd18855: data <= 8'h07;
            16'd18856: data <= 8'hE0;
            16'd18857: data <= 8'h07;
            16'd18858: data <= 8'hE0;
            16'd18859: data <= 8'h07;
            16'd18860: data <= 8'hE0;
            16'd18861: data <= 8'h07;
            16'd18862: data <= 8'hE0;
            16'd18863: data <= 8'h07;
            16'd18864: data <= 8'hE0;
            16'd18865: data <= 8'h07;
            16'd18866: data <= 8'hE0;
            16'd18867: data <= 8'h07;
            16'd18868: data <= 8'hE0;
            16'd18869: data <= 8'h07;
            16'd18870: data <= 8'hE0;
            16'd18871: data <= 8'h07;
            16'd18872: data <= 8'hE0;
            16'd18873: data <= 8'h07;
            16'd18874: data <= 8'hE0;
            16'd18875: data <= 8'h07;
            16'd18876: data <= 8'hE0;
            16'd18877: data <= 8'h07;
            16'd18878: data <= 8'hE0;
            16'd18879: data <= 8'h07;
            16'd18880: data <= 8'hFF;
            16'd18881: data <= 8'hFF;
            16'd18882: data <= 8'hE0;
            16'd18883: data <= 8'h07;
            16'd18884: data <= 8'hE0;
            16'd18885: data <= 8'h07;
            16'd18886: data <= 8'hE0;
            16'd18887: data <= 8'h07;
            16'd18888: data <= 8'hE0;
            16'd18889: data <= 8'h07;
            16'd18890: data <= 8'hE0;
            16'd18891: data <= 8'h07;
            16'd18892: data <= 8'hE0;
            16'd18893: data <= 8'h07;
            16'd18894: data <= 8'hE0;
            16'd18895: data <= 8'h07;
            16'd18896: data <= 8'hE0;
            16'd18897: data <= 8'h07;
            16'd18898: data <= 8'hE0;
            16'd18899: data <= 8'h07;
            16'd18900: data <= 8'hE0;
            16'd18901: data <= 8'h07;
            16'd18902: data <= 8'hE0;
            16'd18903: data <= 8'h07;
            16'd18904: data <= 8'hE0;
            16'd18905: data <= 8'h07;
            16'd18906: data <= 8'hE0;
            16'd18907: data <= 8'h07;
            16'd18908: data <= 8'hE0;
            16'd18909: data <= 8'h07;
            16'd18910: data <= 8'hE0;
            16'd18911: data <= 8'h07;
            16'd18912: data <= 8'hE0;
            16'd18913: data <= 8'h07;
            16'd18914: data <= 8'hE0;
            16'd18915: data <= 8'h07;
            16'd18916: data <= 8'hE0;
            16'd18917: data <= 8'h07;
            16'd18918: data <= 8'hE0;
            16'd18919: data <= 8'h07;
            16'd18920: data <= 8'hFF;
            16'd18921: data <= 8'hFF;
            16'd18922: data <= 8'hE0;
            16'd18923: data <= 8'h07;
            16'd18924: data <= 8'hE0;
            16'd18925: data <= 8'h07;
            16'd18926: data <= 8'hE0;
            16'd18927: data <= 8'h07;
            16'd18928: data <= 8'hE0;
            16'd18929: data <= 8'h07;
            16'd18930: data <= 8'hE0;
            16'd18931: data <= 8'h07;
            16'd18932: data <= 8'hE0;
            16'd18933: data <= 8'h07;
            16'd18934: data <= 8'hE0;
            16'd18935: data <= 8'h07;
            16'd18936: data <= 8'hE0;
            16'd18937: data <= 8'h07;
            16'd18938: data <= 8'hE0;
            16'd18939: data <= 8'h07;
            16'd18940: data <= 8'hE0;
            16'd18941: data <= 8'h07;
            16'd18942: data <= 8'hE0;
            16'd18943: data <= 8'h07;
            16'd18944: data <= 8'hE0;
            16'd18945: data <= 8'h07;
            16'd18946: data <= 8'hE0;
            16'd18947: data <= 8'h07;
            16'd18948: data <= 8'hE0;
            16'd18949: data <= 8'h07;
            16'd18950: data <= 8'hE0;
            16'd18951: data <= 8'h07;
            16'd18952: data <= 8'hE0;
            16'd18953: data <= 8'h07;
            16'd18954: data <= 8'hE0;
            16'd18955: data <= 8'h07;
            16'd18956: data <= 8'hE0;
            16'd18957: data <= 8'h07;
            16'd18958: data <= 8'hE0;
            16'd18959: data <= 8'h07;
            16'd18960: data <= 8'hFF;
            16'd18961: data <= 8'hFF;
            16'd18962: data <= 8'hE0;
            16'd18963: data <= 8'h07;
            16'd18964: data <= 8'hE0;
            16'd18965: data <= 8'h07;
            16'd18966: data <= 8'hE0;
            16'd18967: data <= 8'h07;
            16'd18968: data <= 8'hE0;
            16'd18969: data <= 8'h07;
            16'd18970: data <= 8'hE0;
            16'd18971: data <= 8'h07;
            16'd18972: data <= 8'hE0;
            16'd18973: data <= 8'h07;
            16'd18974: data <= 8'hE0;
            16'd18975: data <= 8'h07;
            16'd18976: data <= 8'hE0;
            16'd18977: data <= 8'h07;
            16'd18978: data <= 8'hE0;
            16'd18979: data <= 8'h07;
            16'd18980: data <= 8'hE0;
            16'd18981: data <= 8'h07;
            16'd18982: data <= 8'hE0;
            16'd18983: data <= 8'h07;
            16'd18984: data <= 8'hE0;
            16'd18985: data <= 8'h07;
            16'd18986: data <= 8'hE0;
            16'd18987: data <= 8'h07;
            16'd18988: data <= 8'hE0;
            16'd18989: data <= 8'h07;
            16'd18990: data <= 8'hE0;
            16'd18991: data <= 8'h07;
            16'd18992: data <= 8'hE0;
            16'd18993: data <= 8'h07;
            16'd18994: data <= 8'hE0;
            16'd18995: data <= 8'h07;
            16'd18996: data <= 8'hE0;
            16'd18997: data <= 8'h07;
            16'd18998: data <= 8'hE0;
            16'd18999: data <= 8'h07;
            16'd19000: data <= 8'hFF;
            16'd19001: data <= 8'hFF;
            16'd19002: data <= 8'hE0;
            16'd19003: data <= 8'h07;
            16'd19004: data <= 8'hE0;
            16'd19005: data <= 8'h07;
            16'd19006: data <= 8'hE0;
            16'd19007: data <= 8'h07;
            16'd19008: data <= 8'hE0;
            16'd19009: data <= 8'h07;
            16'd19010: data <= 8'hE0;
            16'd19011: data <= 8'h07;
            16'd19012: data <= 8'hE0;
            16'd19013: data <= 8'h07;
            16'd19014: data <= 8'hE0;
            16'd19015: data <= 8'h07;
            16'd19016: data <= 8'hE0;
            16'd19017: data <= 8'h07;
            16'd19018: data <= 8'hE0;
            16'd19019: data <= 8'h07;
            16'd19020: data <= 8'hE0;
            16'd19021: data <= 8'h07;
            16'd19022: data <= 8'hE0;
            16'd19023: data <= 8'h07;
            16'd19024: data <= 8'hE0;
            16'd19025: data <= 8'h07;
            16'd19026: data <= 8'hE0;
            16'd19027: data <= 8'h07;
            16'd19028: data <= 8'hE0;
            16'd19029: data <= 8'h07;
            16'd19030: data <= 8'hE0;
            16'd19031: data <= 8'h07;
            16'd19032: data <= 8'hE0;
            16'd19033: data <= 8'h07;
            16'd19034: data <= 8'hE0;
            16'd19035: data <= 8'h07;
            16'd19036: data <= 8'hE0;
            16'd19037: data <= 8'h07;
            16'd19038: data <= 8'hE0;
            16'd19039: data <= 8'h07;
            16'd19040: data <= 8'hFF;
            16'd19041: data <= 8'hFF;
            16'd19042: data <= 8'hE0;
            16'd19043: data <= 8'h07;
            16'd19044: data <= 8'hE0;
            16'd19045: data <= 8'h07;
            16'd19046: data <= 8'hE0;
            16'd19047: data <= 8'h07;
            16'd19048: data <= 8'hE0;
            16'd19049: data <= 8'h07;
            16'd19050: data <= 8'hE0;
            16'd19051: data <= 8'h07;
            16'd19052: data <= 8'hE0;
            16'd19053: data <= 8'h07;
            16'd19054: data <= 8'hE0;
            16'd19055: data <= 8'h07;
            16'd19056: data <= 8'hE0;
            16'd19057: data <= 8'h07;
            16'd19058: data <= 8'hE0;
            16'd19059: data <= 8'h07;
            16'd19060: data <= 8'hE0;
            16'd19061: data <= 8'h07;
            16'd19062: data <= 8'hE0;
            16'd19063: data <= 8'h07;
            16'd19064: data <= 8'hE0;
            16'd19065: data <= 8'h07;
            16'd19066: data <= 8'hE0;
            16'd19067: data <= 8'h07;
            16'd19068: data <= 8'hE0;
            16'd19069: data <= 8'h07;
            16'd19070: data <= 8'hE0;
            16'd19071: data <= 8'h07;
            16'd19072: data <= 8'hE0;
            16'd19073: data <= 8'h07;
            16'd19074: data <= 8'hE0;
            16'd19075: data <= 8'h07;
            16'd19076: data <= 8'hE0;
            16'd19077: data <= 8'h07;
            16'd19078: data <= 8'hE0;
            16'd19079: data <= 8'h07;
            16'd19080: data <= 8'hFF;
            16'd19081: data <= 8'hFF;
            16'd19082: data <= 8'hE0;
            16'd19083: data <= 8'h07;
            16'd19084: data <= 8'hE0;
            16'd19085: data <= 8'h07;
            16'd19086: data <= 8'hE0;
            16'd19087: data <= 8'h07;
            16'd19088: data <= 8'hE0;
            16'd19089: data <= 8'h07;
            16'd19090: data <= 8'hE0;
            16'd19091: data <= 8'h07;
            16'd19092: data <= 8'hE0;
            16'd19093: data <= 8'h07;
            16'd19094: data <= 8'hE0;
            16'd19095: data <= 8'h07;
            16'd19096: data <= 8'hE0;
            16'd19097: data <= 8'h07;
            16'd19098: data <= 8'hE0;
            16'd19099: data <= 8'h07;
            16'd19100: data <= 8'hE0;
            16'd19101: data <= 8'h07;
            16'd19102: data <= 8'hE0;
            16'd19103: data <= 8'h07;
            16'd19104: data <= 8'hE0;
            16'd19105: data <= 8'h07;
            16'd19106: data <= 8'hE0;
            16'd19107: data <= 8'h07;
            16'd19108: data <= 8'hE0;
            16'd19109: data <= 8'h07;
            16'd19110: data <= 8'hE0;
            16'd19111: data <= 8'h07;
            16'd19112: data <= 8'hE0;
            16'd19113: data <= 8'h07;
            16'd19114: data <= 8'hE0;
            16'd19115: data <= 8'h07;
            16'd19116: data <= 8'hE0;
            16'd19117: data <= 8'h07;
            16'd19118: data <= 8'hE0;
            16'd19119: data <= 8'h07;
            16'd19120: data <= 8'hFF;
            16'd19121: data <= 8'hFF;
            16'd19122: data <= 8'hE0;
            16'd19123: data <= 8'h07;
            16'd19124: data <= 8'hE0;
            16'd19125: data <= 8'h07;
            16'd19126: data <= 8'hE0;
            16'd19127: data <= 8'h07;
            16'd19128: data <= 8'hE0;
            16'd19129: data <= 8'h07;
            16'd19130: data <= 8'hE0;
            16'd19131: data <= 8'h07;
            16'd19132: data <= 8'hE0;
            16'd19133: data <= 8'h07;
            16'd19134: data <= 8'hE0;
            16'd19135: data <= 8'h07;
            16'd19136: data <= 8'hE0;
            16'd19137: data <= 8'h07;
            16'd19138: data <= 8'hE0;
            16'd19139: data <= 8'h07;
            16'd19140: data <= 8'hE0;
            16'd19141: data <= 8'h07;
            16'd19142: data <= 8'hE0;
            16'd19143: data <= 8'h07;
            16'd19144: data <= 8'hE0;
            16'd19145: data <= 8'h07;
            16'd19146: data <= 8'hE0;
            16'd19147: data <= 8'h07;
            16'd19148: data <= 8'hE0;
            16'd19149: data <= 8'h07;
            16'd19150: data <= 8'hE0;
            16'd19151: data <= 8'h07;
            16'd19152: data <= 8'hE0;
            16'd19153: data <= 8'h07;
            16'd19154: data <= 8'hE0;
            16'd19155: data <= 8'h07;
            16'd19156: data <= 8'hE0;
            16'd19157: data <= 8'h07;
            16'd19158: data <= 8'hE0;
            16'd19159: data <= 8'h07;
            16'd19160: data <= 8'hFF;
            16'd19161: data <= 8'hFF;
            16'd19162: data <= 8'hE0;
            16'd19163: data <= 8'h07;
            16'd19164: data <= 8'hE0;
            16'd19165: data <= 8'h07;
            16'd19166: data <= 8'hE0;
            16'd19167: data <= 8'h07;
            16'd19168: data <= 8'hE0;
            16'd19169: data <= 8'h07;
            16'd19170: data <= 8'hE0;
            16'd19171: data <= 8'h07;
            16'd19172: data <= 8'hE0;
            16'd19173: data <= 8'h07;
            16'd19174: data <= 8'hE0;
            16'd19175: data <= 8'h07;
            16'd19176: data <= 8'hE0;
            16'd19177: data <= 8'h07;
            16'd19178: data <= 8'hE0;
            16'd19179: data <= 8'h07;
            16'd19180: data <= 8'hE0;
            16'd19181: data <= 8'h07;
            16'd19182: data <= 8'hE0;
            16'd19183: data <= 8'h07;
            16'd19184: data <= 8'hE0;
            16'd19185: data <= 8'h07;
            16'd19186: data <= 8'hE0;
            16'd19187: data <= 8'h07;
            16'd19188: data <= 8'hE0;
            16'd19189: data <= 8'h07;
            16'd19190: data <= 8'hE0;
            16'd19191: data <= 8'h07;
            16'd19192: data <= 8'hE0;
            16'd19193: data <= 8'h07;
            16'd19194: data <= 8'hE0;
            16'd19195: data <= 8'h07;
            16'd19196: data <= 8'hE0;
            16'd19197: data <= 8'h07;
            16'd19198: data <= 8'hE0;
            16'd19199: data <= 8'h07;
            16'd19200: data <= 8'hFF;
            16'd19201: data <= 8'hFF;
            16'd19202: data <= 8'hFF;
            16'd19203: data <= 8'hFF;
            16'd19204: data <= 8'hFF;
            16'd19205: data <= 8'hFF;
            16'd19206: data <= 8'hFF;
            16'd19207: data <= 8'hFF;
            16'd19208: data <= 8'hFF;
            16'd19209: data <= 8'hFF;
            16'd19210: data <= 8'hFF;
            16'd19211: data <= 8'hFF;
            16'd19212: data <= 8'hFF;
            16'd19213: data <= 8'hFF;
            16'd19214: data <= 8'hFF;
            16'd19215: data <= 8'hFF;
            16'd19216: data <= 8'hFF;
            16'd19217: data <= 8'hFF;
            16'd19218: data <= 8'hFF;
            16'd19219: data <= 8'hFF;
            16'd19220: data <= 8'hFF;
            16'd19221: data <= 8'hFF;
            16'd19222: data <= 8'hFF;
            16'd19223: data <= 8'hFF;
            16'd19224: data <= 8'hFF;
            16'd19225: data <= 8'hFF;
            16'd19226: data <= 8'hFF;
            16'd19227: data <= 8'hFF;
            16'd19228: data <= 8'hFF;
            16'd19229: data <= 8'hFF;
            16'd19230: data <= 8'hFF;
            16'd19231: data <= 8'hFF;
            16'd19232: data <= 8'hFF;
            16'd19233: data <= 8'hFF;
            16'd19234: data <= 8'hFF;
            16'd19235: data <= 8'hFF;
            16'd19236: data <= 8'hFF;
            16'd19237: data <= 8'hFF;
            16'd19238: data <= 8'hFF;
            16'd19239: data <= 8'hFF;
            16'd19240: data <= 8'hFF;
            16'd19241: data <= 8'hFF;
            16'd19242: data <= 8'hFF;
            16'd19243: data <= 8'hFF;
            16'd19244: data <= 8'hFF;
            16'd19245: data <= 8'hFF;
            16'd19246: data <= 8'hFF;
            16'd19247: data <= 8'hFF;
            16'd19248: data <= 8'hFF;
            16'd19249: data <= 8'hFF;
            16'd19250: data <= 8'hFF;
            16'd19251: data <= 8'hFF;
            16'd19252: data <= 8'hFF;
            16'd19253: data <= 8'hFF;
            16'd19254: data <= 8'hFF;
            16'd19255: data <= 8'hFF;
            16'd19256: data <= 8'hFF;
            16'd19257: data <= 8'hFF;
            16'd19258: data <= 8'hFF;
            16'd19259: data <= 8'hFF;
            16'd19260: data <= 8'hFF;
            16'd19261: data <= 8'hFF;
            16'd19262: data <= 8'hFF;
            16'd19263: data <= 8'hFF;
            16'd19264: data <= 8'hFF;
            16'd19265: data <= 8'hFF;
            16'd19266: data <= 8'hFF;
            16'd19267: data <= 8'hFF;
            16'd19268: data <= 8'hFF;
            16'd19269: data <= 8'hFF;
            16'd19270: data <= 8'hFF;
            16'd19271: data <= 8'hFF;
            16'd19272: data <= 8'hFF;
            16'd19273: data <= 8'hFF;
            16'd19274: data <= 8'hFF;
            16'd19275: data <= 8'hFF;
            16'd19276: data <= 8'hFF;
            16'd19277: data <= 8'hFF;
            16'd19278: data <= 8'hFF;
            16'd19279: data <= 8'hFF;
            16'd19280: data <= 8'hFF;
            16'd19281: data <= 8'hFF;
            16'd19282: data <= 8'hFF;
            16'd19283: data <= 8'hFF;
            16'd19284: data <= 8'hFF;
            16'd19285: data <= 8'hFF;
            16'd19286: data <= 8'hFF;
            16'd19287: data <= 8'hFF;
            16'd19288: data <= 8'hFF;
            16'd19289: data <= 8'hFF;
            16'd19290: data <= 8'hFF;
            16'd19291: data <= 8'hFF;
            16'd19292: data <= 8'hFF;
            16'd19293: data <= 8'hFF;
            16'd19294: data <= 8'hFF;
            16'd19295: data <= 8'hFF;
            16'd19296: data <= 8'hFF;
            16'd19297: data <= 8'hFF;
            16'd19298: data <= 8'hFF;
            16'd19299: data <= 8'hFF;
            16'd19300: data <= 8'hFF;
            16'd19301: data <= 8'hFF;
            16'd19302: data <= 8'hFF;
            16'd19303: data <= 8'hFF;
            16'd19304: data <= 8'hFF;
            16'd19305: data <= 8'hFF;
            16'd19306: data <= 8'hFF;
            16'd19307: data <= 8'hFF;
            16'd19308: data <= 8'hFF;
            16'd19309: data <= 8'hFF;
            16'd19310: data <= 8'hFF;
            16'd19311: data <= 8'hFF;
            16'd19312: data <= 8'hFF;
            16'd19313: data <= 8'hFF;
            16'd19314: data <= 8'hFF;
            16'd19315: data <= 8'hFF;
            16'd19316: data <= 8'hFF;
            16'd19317: data <= 8'hFF;
            16'd19318: data <= 8'hFF;
            16'd19319: data <= 8'hFF;
            16'd19320: data <= 8'hFF;
            16'd19321: data <= 8'hFF;
            16'd19322: data <= 8'hFF;
            16'd19323: data <= 8'hFF;
            16'd19324: data <= 8'hFF;
            16'd19325: data <= 8'hFF;
            16'd19326: data <= 8'hFF;
            16'd19327: data <= 8'hFF;
            16'd19328: data <= 8'hFF;
            16'd19329: data <= 8'hFF;
            16'd19330: data <= 8'hFF;
            16'd19331: data <= 8'hFF;
            16'd19332: data <= 8'hFF;
            16'd19333: data <= 8'hFF;
            16'd19334: data <= 8'hFF;
            16'd19335: data <= 8'hFF;
            16'd19336: data <= 8'hFF;
            16'd19337: data <= 8'hFF;
            16'd19338: data <= 8'hFF;
            16'd19339: data <= 8'hFF;
            16'd19340: data <= 8'hFF;
            16'd19341: data <= 8'hFF;
            16'd19342: data <= 8'hFF;
            16'd19343: data <= 8'hFF;
            16'd19344: data <= 8'hFF;
            16'd19345: data <= 8'hFF;
            16'd19346: data <= 8'hFF;
            16'd19347: data <= 8'hFF;
            16'd19348: data <= 8'hFF;
            16'd19349: data <= 8'hFF;
            16'd19350: data <= 8'hFF;
            16'd19351: data <= 8'hFF;
            16'd19352: data <= 8'hFF;
            16'd19353: data <= 8'hFF;
            16'd19354: data <= 8'hFF;
            16'd19355: data <= 8'hFF;
            16'd19356: data <= 8'hFF;
            16'd19357: data <= 8'hFF;
            16'd19358: data <= 8'hFF;
            16'd19359: data <= 8'hFF;
            16'd19360: data <= 8'hFF;
            16'd19361: data <= 8'hFF;
            16'd19362: data <= 8'hFF;
            16'd19363: data <= 8'hFF;
            16'd19364: data <= 8'hFF;
            16'd19365: data <= 8'hFF;
            16'd19366: data <= 8'hFF;
            16'd19367: data <= 8'hFF;
            16'd19368: data <= 8'hFF;
            16'd19369: data <= 8'hFF;
            16'd19370: data <= 8'hFF;
            16'd19371: data <= 8'hFF;
            16'd19372: data <= 8'hFF;
            16'd19373: data <= 8'hFF;
            16'd19374: data <= 8'hFF;
            16'd19375: data <= 8'hFF;
            16'd19376: data <= 8'hFF;
            16'd19377: data <= 8'hFF;
            16'd19378: data <= 8'hFF;
            16'd19379: data <= 8'hFF;
            16'd19380: data <= 8'hFF;
            16'd19381: data <= 8'hFF;
            16'd19382: data <= 8'hFF;
            16'd19383: data <= 8'hFF;
            16'd19384: data <= 8'hFF;
            16'd19385: data <= 8'hFF;
            16'd19386: data <= 8'hFF;
            16'd19387: data <= 8'hFF;
            16'd19388: data <= 8'hFF;
            16'd19389: data <= 8'hFF;
            16'd19390: data <= 8'hFF;
            16'd19391: data <= 8'hFF;
            16'd19392: data <= 8'hFF;
            16'd19393: data <= 8'hFF;
            16'd19394: data <= 8'hFF;
            16'd19395: data <= 8'hFF;
            16'd19396: data <= 8'hFF;
            16'd19397: data <= 8'hFF;
            16'd19398: data <= 8'hFF;
            16'd19399: data <= 8'hFF;
            16'd19400: data <= 8'hFF;
            16'd19401: data <= 8'hFF;
            16'd19402: data <= 8'hFF;
            16'd19403: data <= 8'hFF;
            16'd19404: data <= 8'hFF;
            16'd19405: data <= 8'hFF;
            16'd19406: data <= 8'hFF;
            16'd19407: data <= 8'hFF;
            16'd19408: data <= 8'hFF;
            16'd19409: data <= 8'hFF;
            16'd19410: data <= 8'hFF;
            16'd19411: data <= 8'hFF;
            16'd19412: data <= 8'hFF;
            16'd19413: data <= 8'hFF;
            16'd19414: data <= 8'hFF;
            16'd19415: data <= 8'hFF;
            16'd19416: data <= 8'hFF;
            16'd19417: data <= 8'hFF;
            16'd19418: data <= 8'hFF;
            16'd19419: data <= 8'hFF;
            16'd19420: data <= 8'hFF;
            16'd19421: data <= 8'hFF;
            16'd19422: data <= 8'hFF;
            16'd19423: data <= 8'hFF;
            16'd19424: data <= 8'hFF;
            16'd19425: data <= 8'hFF;
            16'd19426: data <= 8'hFF;
            16'd19427: data <= 8'hFF;
            16'd19428: data <= 8'hFF;
            16'd19429: data <= 8'hFF;
            16'd19430: data <= 8'hFF;
            16'd19431: data <= 8'hFF;
            16'd19432: data <= 8'hFF;
            16'd19433: data <= 8'hFF;
            16'd19434: data <= 8'hFF;
            16'd19435: data <= 8'hFF;
            16'd19436: data <= 8'hFF;
            16'd19437: data <= 8'hFF;
            16'd19438: data <= 8'hFF;
            16'd19439: data <= 8'hFF;
            16'd19440: data <= 8'hFF;
            16'd19441: data <= 8'hFF;
            16'd19442: data <= 8'hE0;
            16'd19443: data <= 8'h07;
            16'd19444: data <= 8'hE0;
            16'd19445: data <= 8'h07;
            16'd19446: data <= 8'hE0;
            16'd19447: data <= 8'h07;
            16'd19448: data <= 8'hE0;
            16'd19449: data <= 8'h07;
            16'd19450: data <= 8'hE0;
            16'd19451: data <= 8'h07;
            16'd19452: data <= 8'hE0;
            16'd19453: data <= 8'h07;
            16'd19454: data <= 8'hE0;
            16'd19455: data <= 8'h07;
            16'd19456: data <= 8'hE0;
            16'd19457: data <= 8'h07;
            16'd19458: data <= 8'hE0;
            16'd19459: data <= 8'h07;
            16'd19460: data <= 8'hE0;
            16'd19461: data <= 8'h07;
            16'd19462: data <= 8'hE0;
            16'd19463: data <= 8'h07;
            16'd19464: data <= 8'hE0;
            16'd19465: data <= 8'h07;
            16'd19466: data <= 8'hE0;
            16'd19467: data <= 8'h07;
            16'd19468: data <= 8'hE0;
            16'd19469: data <= 8'h07;
            16'd19470: data <= 8'hE0;
            16'd19471: data <= 8'h07;
            16'd19472: data <= 8'hE0;
            16'd19473: data <= 8'h07;
            16'd19474: data <= 8'hE0;
            16'd19475: data <= 8'h07;
            16'd19476: data <= 8'hE0;
            16'd19477: data <= 8'h07;
            16'd19478: data <= 8'hE0;
            16'd19479: data <= 8'h07;
            16'd19480: data <= 8'hFF;
            16'd19481: data <= 8'hFF;
            16'd19482: data <= 8'hE0;
            16'd19483: data <= 8'h07;
            16'd19484: data <= 8'hE0;
            16'd19485: data <= 8'h07;
            16'd19486: data <= 8'hE0;
            16'd19487: data <= 8'h07;
            16'd19488: data <= 8'hE0;
            16'd19489: data <= 8'h07;
            16'd19490: data <= 8'hE0;
            16'd19491: data <= 8'h07;
            16'd19492: data <= 8'hE0;
            16'd19493: data <= 8'h07;
            16'd19494: data <= 8'hE0;
            16'd19495: data <= 8'h07;
            16'd19496: data <= 8'hE0;
            16'd19497: data <= 8'h07;
            16'd19498: data <= 8'hE0;
            16'd19499: data <= 8'h07;
            16'd19500: data <= 8'hE0;
            16'd19501: data <= 8'h07;
            16'd19502: data <= 8'hE0;
            16'd19503: data <= 8'h07;
            16'd19504: data <= 8'hE0;
            16'd19505: data <= 8'h07;
            16'd19506: data <= 8'hE0;
            16'd19507: data <= 8'h07;
            16'd19508: data <= 8'hE0;
            16'd19509: data <= 8'h07;
            16'd19510: data <= 8'hE0;
            16'd19511: data <= 8'h07;
            16'd19512: data <= 8'hE0;
            16'd19513: data <= 8'h07;
            16'd19514: data <= 8'hE0;
            16'd19515: data <= 8'h07;
            16'd19516: data <= 8'hE0;
            16'd19517: data <= 8'h07;
            16'd19518: data <= 8'hE0;
            16'd19519: data <= 8'h07;
            16'd19520: data <= 8'hFF;
            16'd19521: data <= 8'hFF;
            16'd19522: data <= 8'hE0;
            16'd19523: data <= 8'h07;
            16'd19524: data <= 8'hE0;
            16'd19525: data <= 8'h07;
            16'd19526: data <= 8'hE0;
            16'd19527: data <= 8'h07;
            16'd19528: data <= 8'hE0;
            16'd19529: data <= 8'h07;
            16'd19530: data <= 8'hE0;
            16'd19531: data <= 8'h07;
            16'd19532: data <= 8'hE0;
            16'd19533: data <= 8'h07;
            16'd19534: data <= 8'hE0;
            16'd19535: data <= 8'h07;
            16'd19536: data <= 8'hE0;
            16'd19537: data <= 8'h07;
            16'd19538: data <= 8'hE0;
            16'd19539: data <= 8'h07;
            16'd19540: data <= 8'hE0;
            16'd19541: data <= 8'h07;
            16'd19542: data <= 8'hE0;
            16'd19543: data <= 8'h07;
            16'd19544: data <= 8'hE0;
            16'd19545: data <= 8'h07;
            16'd19546: data <= 8'hE0;
            16'd19547: data <= 8'h07;
            16'd19548: data <= 8'hE0;
            16'd19549: data <= 8'h07;
            16'd19550: data <= 8'hE0;
            16'd19551: data <= 8'h07;
            16'd19552: data <= 8'hE0;
            16'd19553: data <= 8'h07;
            16'd19554: data <= 8'hE0;
            16'd19555: data <= 8'h07;
            16'd19556: data <= 8'hE0;
            16'd19557: data <= 8'h07;
            16'd19558: data <= 8'hE0;
            16'd19559: data <= 8'h07;
            16'd19560: data <= 8'hFF;
            16'd19561: data <= 8'hFF;
            16'd19562: data <= 8'hE0;
            16'd19563: data <= 8'h07;
            16'd19564: data <= 8'hE0;
            16'd19565: data <= 8'h07;
            16'd19566: data <= 8'hE0;
            16'd19567: data <= 8'h07;
            16'd19568: data <= 8'hE0;
            16'd19569: data <= 8'h07;
            16'd19570: data <= 8'hE0;
            16'd19571: data <= 8'h07;
            16'd19572: data <= 8'hE0;
            16'd19573: data <= 8'h07;
            16'd19574: data <= 8'hE0;
            16'd19575: data <= 8'h07;
            16'd19576: data <= 8'hE0;
            16'd19577: data <= 8'h07;
            16'd19578: data <= 8'hE0;
            16'd19579: data <= 8'h07;
            16'd19580: data <= 8'hE0;
            16'd19581: data <= 8'h07;
            16'd19582: data <= 8'hE0;
            16'd19583: data <= 8'h07;
            16'd19584: data <= 8'hE0;
            16'd19585: data <= 8'h07;
            16'd19586: data <= 8'hE0;
            16'd19587: data <= 8'h07;
            16'd19588: data <= 8'hE0;
            16'd19589: data <= 8'h07;
            16'd19590: data <= 8'hE0;
            16'd19591: data <= 8'h07;
            16'd19592: data <= 8'hE0;
            16'd19593: data <= 8'h07;
            16'd19594: data <= 8'hE0;
            16'd19595: data <= 8'h07;
            16'd19596: data <= 8'hE0;
            16'd19597: data <= 8'h07;
            16'd19598: data <= 8'hE0;
            16'd19599: data <= 8'h07;
            16'd19600: data <= 8'hFF;
            16'd19601: data <= 8'hFF;
            16'd19602: data <= 8'hE0;
            16'd19603: data <= 8'h07;
            16'd19604: data <= 8'hE0;
            16'd19605: data <= 8'h07;
            16'd19606: data <= 8'hE0;
            16'd19607: data <= 8'h07;
            16'd19608: data <= 8'hE0;
            16'd19609: data <= 8'h07;
            16'd19610: data <= 8'hE0;
            16'd19611: data <= 8'h07;
            16'd19612: data <= 8'hE0;
            16'd19613: data <= 8'h07;
            16'd19614: data <= 8'hE0;
            16'd19615: data <= 8'h07;
            16'd19616: data <= 8'hE0;
            16'd19617: data <= 8'h07;
            16'd19618: data <= 8'hE0;
            16'd19619: data <= 8'h07;
            16'd19620: data <= 8'hE0;
            16'd19621: data <= 8'h07;
            16'd19622: data <= 8'hE0;
            16'd19623: data <= 8'h07;
            16'd19624: data <= 8'hE0;
            16'd19625: data <= 8'h07;
            16'd19626: data <= 8'hE0;
            16'd19627: data <= 8'h07;
            16'd19628: data <= 8'hE0;
            16'd19629: data <= 8'h07;
            16'd19630: data <= 8'hE0;
            16'd19631: data <= 8'h07;
            16'd19632: data <= 8'hE0;
            16'd19633: data <= 8'h07;
            16'd19634: data <= 8'hE0;
            16'd19635: data <= 8'h07;
            16'd19636: data <= 8'hE0;
            16'd19637: data <= 8'h07;
            16'd19638: data <= 8'hE0;
            16'd19639: data <= 8'h07;
            16'd19640: data <= 8'hFF;
            16'd19641: data <= 8'hFF;
            16'd19642: data <= 8'hE0;
            16'd19643: data <= 8'h07;
            16'd19644: data <= 8'hE0;
            16'd19645: data <= 8'h07;
            16'd19646: data <= 8'hE0;
            16'd19647: data <= 8'h07;
            16'd19648: data <= 8'hE0;
            16'd19649: data <= 8'h07;
            16'd19650: data <= 8'hE0;
            16'd19651: data <= 8'h07;
            16'd19652: data <= 8'hE0;
            16'd19653: data <= 8'h07;
            16'd19654: data <= 8'hE0;
            16'd19655: data <= 8'h07;
            16'd19656: data <= 8'hE0;
            16'd19657: data <= 8'h07;
            16'd19658: data <= 8'hE0;
            16'd19659: data <= 8'h07;
            16'd19660: data <= 8'hE0;
            16'd19661: data <= 8'h07;
            16'd19662: data <= 8'hE0;
            16'd19663: data <= 8'h07;
            16'd19664: data <= 8'hE0;
            16'd19665: data <= 8'h07;
            16'd19666: data <= 8'hE0;
            16'd19667: data <= 8'h07;
            16'd19668: data <= 8'hE0;
            16'd19669: data <= 8'h07;
            16'd19670: data <= 8'hE0;
            16'd19671: data <= 8'h07;
            16'd19672: data <= 8'hE0;
            16'd19673: data <= 8'h07;
            16'd19674: data <= 8'hE0;
            16'd19675: data <= 8'h07;
            16'd19676: data <= 8'hE0;
            16'd19677: data <= 8'h07;
            16'd19678: data <= 8'hE0;
            16'd19679: data <= 8'h07;
            16'd19680: data <= 8'hFF;
            16'd19681: data <= 8'hFF;
            16'd19682: data <= 8'hE0;
            16'd19683: data <= 8'h07;
            16'd19684: data <= 8'hE0;
            16'd19685: data <= 8'h07;
            16'd19686: data <= 8'hE0;
            16'd19687: data <= 8'h07;
            16'd19688: data <= 8'hE0;
            16'd19689: data <= 8'h07;
            16'd19690: data <= 8'hE0;
            16'd19691: data <= 8'h07;
            16'd19692: data <= 8'hE0;
            16'd19693: data <= 8'h07;
            16'd19694: data <= 8'hE0;
            16'd19695: data <= 8'h07;
            16'd19696: data <= 8'hE0;
            16'd19697: data <= 8'h07;
            16'd19698: data <= 8'hE0;
            16'd19699: data <= 8'h07;
            16'd19700: data <= 8'hE0;
            16'd19701: data <= 8'h07;
            16'd19702: data <= 8'hE0;
            16'd19703: data <= 8'h07;
            16'd19704: data <= 8'hE0;
            16'd19705: data <= 8'h07;
            16'd19706: data <= 8'hE0;
            16'd19707: data <= 8'h07;
            16'd19708: data <= 8'hE0;
            16'd19709: data <= 8'h07;
            16'd19710: data <= 8'hE0;
            16'd19711: data <= 8'h07;
            16'd19712: data <= 8'hE0;
            16'd19713: data <= 8'h07;
            16'd19714: data <= 8'hE0;
            16'd19715: data <= 8'h07;
            16'd19716: data <= 8'hE0;
            16'd19717: data <= 8'h07;
            16'd19718: data <= 8'hE0;
            16'd19719: data <= 8'h07;
            16'd19720: data <= 8'hFF;
            16'd19721: data <= 8'hFF;
            16'd19722: data <= 8'hE0;
            16'd19723: data <= 8'h07;
            16'd19724: data <= 8'hE0;
            16'd19725: data <= 8'h07;
            16'd19726: data <= 8'hE0;
            16'd19727: data <= 8'h07;
            16'd19728: data <= 8'hE0;
            16'd19729: data <= 8'h07;
            16'd19730: data <= 8'hE0;
            16'd19731: data <= 8'h07;
            16'd19732: data <= 8'hE0;
            16'd19733: data <= 8'h07;
            16'd19734: data <= 8'hE0;
            16'd19735: data <= 8'h07;
            16'd19736: data <= 8'hE0;
            16'd19737: data <= 8'h07;
            16'd19738: data <= 8'hE0;
            16'd19739: data <= 8'h07;
            16'd19740: data <= 8'hE0;
            16'd19741: data <= 8'h07;
            16'd19742: data <= 8'hE0;
            16'd19743: data <= 8'h07;
            16'd19744: data <= 8'hE0;
            16'd19745: data <= 8'h07;
            16'd19746: data <= 8'hE0;
            16'd19747: data <= 8'h07;
            16'd19748: data <= 8'hE0;
            16'd19749: data <= 8'h07;
            16'd19750: data <= 8'hE0;
            16'd19751: data <= 8'h07;
            16'd19752: data <= 8'hE0;
            16'd19753: data <= 8'h07;
            16'd19754: data <= 8'hE0;
            16'd19755: data <= 8'h07;
            16'd19756: data <= 8'hE0;
            16'd19757: data <= 8'h07;
            16'd19758: data <= 8'hE0;
            16'd19759: data <= 8'h07;
            16'd19760: data <= 8'hFF;
            16'd19761: data <= 8'hFF;
            16'd19762: data <= 8'hE0;
            16'd19763: data <= 8'h07;
            16'd19764: data <= 8'hE0;
            16'd19765: data <= 8'h07;
            16'd19766: data <= 8'hE0;
            16'd19767: data <= 8'h07;
            16'd19768: data <= 8'hE0;
            16'd19769: data <= 8'h07;
            16'd19770: data <= 8'hE0;
            16'd19771: data <= 8'h07;
            16'd19772: data <= 8'hE0;
            16'd19773: data <= 8'h07;
            16'd19774: data <= 8'hE0;
            16'd19775: data <= 8'h07;
            16'd19776: data <= 8'hE0;
            16'd19777: data <= 8'h07;
            16'd19778: data <= 8'hE0;
            16'd19779: data <= 8'h07;
            16'd19780: data <= 8'hE0;
            16'd19781: data <= 8'h07;
            16'd19782: data <= 8'hE0;
            16'd19783: data <= 8'h07;
            16'd19784: data <= 8'hE0;
            16'd19785: data <= 8'h07;
            16'd19786: data <= 8'hE0;
            16'd19787: data <= 8'h07;
            16'd19788: data <= 8'hE0;
            16'd19789: data <= 8'h07;
            16'd19790: data <= 8'hE0;
            16'd19791: data <= 8'h07;
            16'd19792: data <= 8'hE0;
            16'd19793: data <= 8'h07;
            16'd19794: data <= 8'hE0;
            16'd19795: data <= 8'h07;
            16'd19796: data <= 8'hE0;
            16'd19797: data <= 8'h07;
            16'd19798: data <= 8'hE0;
            16'd19799: data <= 8'h07;
            16'd19800: data <= 8'hFF;
            16'd19801: data <= 8'hFF;
            16'd19802: data <= 8'hE0;
            16'd19803: data <= 8'h07;
            16'd19804: data <= 8'hE0;
            16'd19805: data <= 8'h07;
            16'd19806: data <= 8'hE0;
            16'd19807: data <= 8'h07;
            16'd19808: data <= 8'hE0;
            16'd19809: data <= 8'h07;
            16'd19810: data <= 8'hE0;
            16'd19811: data <= 8'h07;
            16'd19812: data <= 8'hE0;
            16'd19813: data <= 8'h07;
            16'd19814: data <= 8'hE0;
            16'd19815: data <= 8'h07;
            16'd19816: data <= 8'hE0;
            16'd19817: data <= 8'h07;
            16'd19818: data <= 8'hE0;
            16'd19819: data <= 8'h07;
            16'd19820: data <= 8'hE0;
            16'd19821: data <= 8'h07;
            16'd19822: data <= 8'hE0;
            16'd19823: data <= 8'h07;
            16'd19824: data <= 8'hE0;
            16'd19825: data <= 8'h07;
            16'd19826: data <= 8'hE0;
            16'd19827: data <= 8'h07;
            16'd19828: data <= 8'hE0;
            16'd19829: data <= 8'h07;
            16'd19830: data <= 8'hE0;
            16'd19831: data <= 8'h07;
            16'd19832: data <= 8'hE0;
            16'd19833: data <= 8'h07;
            16'd19834: data <= 8'hE0;
            16'd19835: data <= 8'h07;
            16'd19836: data <= 8'hE0;
            16'd19837: data <= 8'h07;
            16'd19838: data <= 8'hE0;
            16'd19839: data <= 8'h07;
            16'd19840: data <= 8'hFF;
            16'd19841: data <= 8'hFF;
            16'd19842: data <= 8'hE0;
            16'd19843: data <= 8'h07;
            16'd19844: data <= 8'hE0;
            16'd19845: data <= 8'h07;
            16'd19846: data <= 8'hE0;
            16'd19847: data <= 8'h07;
            16'd19848: data <= 8'hE0;
            16'd19849: data <= 8'h07;
            16'd19850: data <= 8'hE0;
            16'd19851: data <= 8'h07;
            16'd19852: data <= 8'hE0;
            16'd19853: data <= 8'h07;
            16'd19854: data <= 8'hE0;
            16'd19855: data <= 8'h07;
            16'd19856: data <= 8'hE0;
            16'd19857: data <= 8'h07;
            16'd19858: data <= 8'hE0;
            16'd19859: data <= 8'h07;
            16'd19860: data <= 8'hE0;
            16'd19861: data <= 8'h07;
            16'd19862: data <= 8'hE0;
            16'd19863: data <= 8'h07;
            16'd19864: data <= 8'hE0;
            16'd19865: data <= 8'h07;
            16'd19866: data <= 8'hE0;
            16'd19867: data <= 8'h07;
            16'd19868: data <= 8'hE0;
            16'd19869: data <= 8'h07;
            16'd19870: data <= 8'hE0;
            16'd19871: data <= 8'h07;
            16'd19872: data <= 8'hE0;
            16'd19873: data <= 8'h07;
            16'd19874: data <= 8'hE0;
            16'd19875: data <= 8'h07;
            16'd19876: data <= 8'hE0;
            16'd19877: data <= 8'h07;
            16'd19878: data <= 8'hE0;
            16'd19879: data <= 8'h07;
            16'd19880: data <= 8'hFF;
            16'd19881: data <= 8'hFF;
            16'd19882: data <= 8'hE0;
            16'd19883: data <= 8'h07;
            16'd19884: data <= 8'hE0;
            16'd19885: data <= 8'h07;
            16'd19886: data <= 8'hE0;
            16'd19887: data <= 8'h07;
            16'd19888: data <= 8'hE0;
            16'd19889: data <= 8'h07;
            16'd19890: data <= 8'hE0;
            16'd19891: data <= 8'h07;
            16'd19892: data <= 8'hE0;
            16'd19893: data <= 8'h07;
            16'd19894: data <= 8'hE0;
            16'd19895: data <= 8'h07;
            16'd19896: data <= 8'hE0;
            16'd19897: data <= 8'h07;
            16'd19898: data <= 8'hE0;
            16'd19899: data <= 8'h07;
            16'd19900: data <= 8'hE0;
            16'd19901: data <= 8'h07;
            16'd19902: data <= 8'hE0;
            16'd19903: data <= 8'h07;
            16'd19904: data <= 8'hE0;
            16'd19905: data <= 8'h07;
            16'd19906: data <= 8'hE0;
            16'd19907: data <= 8'h07;
            16'd19908: data <= 8'hE0;
            16'd19909: data <= 8'h07;
            16'd19910: data <= 8'hE0;
            16'd19911: data <= 8'h07;
            16'd19912: data <= 8'hE0;
            16'd19913: data <= 8'h07;
            16'd19914: data <= 8'hE0;
            16'd19915: data <= 8'h07;
            16'd19916: data <= 8'hE0;
            16'd19917: data <= 8'h07;
            16'd19918: data <= 8'hE0;
            16'd19919: data <= 8'h07;
            16'd19920: data <= 8'hFF;
            16'd19921: data <= 8'hFF;
            16'd19922: data <= 8'hE0;
            16'd19923: data <= 8'h07;
            16'd19924: data <= 8'hE0;
            16'd19925: data <= 8'h07;
            16'd19926: data <= 8'hE0;
            16'd19927: data <= 8'h07;
            16'd19928: data <= 8'hE0;
            16'd19929: data <= 8'h07;
            16'd19930: data <= 8'hE0;
            16'd19931: data <= 8'h07;
            16'd19932: data <= 8'hE0;
            16'd19933: data <= 8'h07;
            16'd19934: data <= 8'hE0;
            16'd19935: data <= 8'h07;
            16'd19936: data <= 8'hE0;
            16'd19937: data <= 8'h07;
            16'd19938: data <= 8'hE0;
            16'd19939: data <= 8'h07;
            16'd19940: data <= 8'hE0;
            16'd19941: data <= 8'h07;
            16'd19942: data <= 8'hE0;
            16'd19943: data <= 8'h07;
            16'd19944: data <= 8'hE0;
            16'd19945: data <= 8'h07;
            16'd19946: data <= 8'hE0;
            16'd19947: data <= 8'h07;
            16'd19948: data <= 8'hE0;
            16'd19949: data <= 8'h07;
            16'd19950: data <= 8'hE0;
            16'd19951: data <= 8'h07;
            16'd19952: data <= 8'hE0;
            16'd19953: data <= 8'h07;
            16'd19954: data <= 8'hE0;
            16'd19955: data <= 8'h07;
            16'd19956: data <= 8'hE0;
            16'd19957: data <= 8'h07;
            16'd19958: data <= 8'hE0;
            16'd19959: data <= 8'h07;
            16'd19960: data <= 8'hFF;
            16'd19961: data <= 8'hFF;
            16'd19962: data <= 8'hE0;
            16'd19963: data <= 8'h07;
            16'd19964: data <= 8'hE0;
            16'd19965: data <= 8'h07;
            16'd19966: data <= 8'hE0;
            16'd19967: data <= 8'h07;
            16'd19968: data <= 8'hE0;
            16'd19969: data <= 8'h07;
            16'd19970: data <= 8'hE0;
            16'd19971: data <= 8'h07;
            16'd19972: data <= 8'hE0;
            16'd19973: data <= 8'h07;
            16'd19974: data <= 8'hE0;
            16'd19975: data <= 8'h07;
            16'd19976: data <= 8'hE0;
            16'd19977: data <= 8'h07;
            16'd19978: data <= 8'hE0;
            16'd19979: data <= 8'h07;
            16'd19980: data <= 8'hE0;
            16'd19981: data <= 8'h07;
            16'd19982: data <= 8'hE0;
            16'd19983: data <= 8'h07;
            16'd19984: data <= 8'hE0;
            16'd19985: data <= 8'h07;
            16'd19986: data <= 8'hE0;
            16'd19987: data <= 8'h07;
            16'd19988: data <= 8'hE0;
            16'd19989: data <= 8'h07;
            16'd19990: data <= 8'hE0;
            16'd19991: data <= 8'h07;
            16'd19992: data <= 8'hE0;
            16'd19993: data <= 8'h07;
            16'd19994: data <= 8'hE0;
            16'd19995: data <= 8'h07;
            16'd19996: data <= 8'hE0;
            16'd19997: data <= 8'h07;
            16'd19998: data <= 8'hE0;
            16'd19999: data <= 8'h07;
            16'd20000: data <= 8'hFF;
            16'd20001: data <= 8'hFF;
            16'd20002: data <= 8'hE0;
            16'd20003: data <= 8'h07;
            16'd20004: data <= 8'hE0;
            16'd20005: data <= 8'h07;
            16'd20006: data <= 8'hE0;
            16'd20007: data <= 8'h07;
            16'd20008: data <= 8'hE0;
            16'd20009: data <= 8'h07;
            16'd20010: data <= 8'hE0;
            16'd20011: data <= 8'h07;
            16'd20012: data <= 8'hE0;
            16'd20013: data <= 8'h07;
            16'd20014: data <= 8'hE0;
            16'd20015: data <= 8'h07;
            16'd20016: data <= 8'hE0;
            16'd20017: data <= 8'h07;
            16'd20018: data <= 8'hE0;
            16'd20019: data <= 8'h07;
            16'd20020: data <= 8'hE0;
            16'd20021: data <= 8'h07;
            16'd20022: data <= 8'hE0;
            16'd20023: data <= 8'h07;
            16'd20024: data <= 8'hE0;
            16'd20025: data <= 8'h07;
            16'd20026: data <= 8'hE0;
            16'd20027: data <= 8'h07;
            16'd20028: data <= 8'hE0;
            16'd20029: data <= 8'h07;
            16'd20030: data <= 8'hE0;
            16'd20031: data <= 8'h07;
            16'd20032: data <= 8'hE0;
            16'd20033: data <= 8'h07;
            16'd20034: data <= 8'hE0;
            16'd20035: data <= 8'h07;
            16'd20036: data <= 8'hE0;
            16'd20037: data <= 8'h07;
            16'd20038: data <= 8'hE0;
            16'd20039: data <= 8'h07;
            16'd20040: data <= 8'hFF;
            16'd20041: data <= 8'hFF;
            16'd20042: data <= 8'hE0;
            16'd20043: data <= 8'h07;
            16'd20044: data <= 8'hE0;
            16'd20045: data <= 8'h07;
            16'd20046: data <= 8'hE0;
            16'd20047: data <= 8'h07;
            16'd20048: data <= 8'hE0;
            16'd20049: data <= 8'h07;
            16'd20050: data <= 8'hE0;
            16'd20051: data <= 8'h07;
            16'd20052: data <= 8'hE0;
            16'd20053: data <= 8'h07;
            16'd20054: data <= 8'hE0;
            16'd20055: data <= 8'h07;
            16'd20056: data <= 8'hE0;
            16'd20057: data <= 8'h07;
            16'd20058: data <= 8'hE0;
            16'd20059: data <= 8'h07;
            16'd20060: data <= 8'hE0;
            16'd20061: data <= 8'h07;
            16'd20062: data <= 8'hE0;
            16'd20063: data <= 8'h07;
            16'd20064: data <= 8'hE0;
            16'd20065: data <= 8'h07;
            16'd20066: data <= 8'hE0;
            16'd20067: data <= 8'h07;
            16'd20068: data <= 8'hE0;
            16'd20069: data <= 8'h07;
            16'd20070: data <= 8'hE0;
            16'd20071: data <= 8'h07;
            16'd20072: data <= 8'hE0;
            16'd20073: data <= 8'h07;
            16'd20074: data <= 8'hE0;
            16'd20075: data <= 8'h07;
            16'd20076: data <= 8'hE0;
            16'd20077: data <= 8'h07;
            16'd20078: data <= 8'hE0;
            16'd20079: data <= 8'h07;
            16'd20080: data <= 8'hFF;
            16'd20081: data <= 8'hFF;
            16'd20082: data <= 8'hE0;
            16'd20083: data <= 8'h07;
            16'd20084: data <= 8'hE0;
            16'd20085: data <= 8'h07;
            16'd20086: data <= 8'hE0;
            16'd20087: data <= 8'h07;
            16'd20088: data <= 8'hE0;
            16'd20089: data <= 8'h07;
            16'd20090: data <= 8'hE0;
            16'd20091: data <= 8'h07;
            16'd20092: data <= 8'hE0;
            16'd20093: data <= 8'h07;
            16'd20094: data <= 8'hE0;
            16'd20095: data <= 8'h07;
            16'd20096: data <= 8'hE0;
            16'd20097: data <= 8'h07;
            16'd20098: data <= 8'hE0;
            16'd20099: data <= 8'h07;
            16'd20100: data <= 8'hE0;
            16'd20101: data <= 8'h07;
            16'd20102: data <= 8'hE0;
            16'd20103: data <= 8'h07;
            16'd20104: data <= 8'hE0;
            16'd20105: data <= 8'h07;
            16'd20106: data <= 8'hE0;
            16'd20107: data <= 8'h07;
            16'd20108: data <= 8'hE0;
            16'd20109: data <= 8'h07;
            16'd20110: data <= 8'hE0;
            16'd20111: data <= 8'h07;
            16'd20112: data <= 8'hE0;
            16'd20113: data <= 8'h07;
            16'd20114: data <= 8'hE0;
            16'd20115: data <= 8'h07;
            16'd20116: data <= 8'hE0;
            16'd20117: data <= 8'h07;
            16'd20118: data <= 8'hE0;
            16'd20119: data <= 8'h07;
            16'd20120: data <= 8'hFF;
            16'd20121: data <= 8'hFF;
            16'd20122: data <= 8'hE0;
            16'd20123: data <= 8'h07;
            16'd20124: data <= 8'hE0;
            16'd20125: data <= 8'h07;
            16'd20126: data <= 8'hE0;
            16'd20127: data <= 8'h07;
            16'd20128: data <= 8'hE0;
            16'd20129: data <= 8'h07;
            16'd20130: data <= 8'hE0;
            16'd20131: data <= 8'h07;
            16'd20132: data <= 8'hE0;
            16'd20133: data <= 8'h07;
            16'd20134: data <= 8'hE0;
            16'd20135: data <= 8'h07;
            16'd20136: data <= 8'hE0;
            16'd20137: data <= 8'h07;
            16'd20138: data <= 8'hE0;
            16'd20139: data <= 8'h07;
            16'd20140: data <= 8'hE0;
            16'd20141: data <= 8'h07;
            16'd20142: data <= 8'hE0;
            16'd20143: data <= 8'h07;
            16'd20144: data <= 8'hE0;
            16'd20145: data <= 8'h07;
            16'd20146: data <= 8'hE0;
            16'd20147: data <= 8'h07;
            16'd20148: data <= 8'hE0;
            16'd20149: data <= 8'h07;
            16'd20150: data <= 8'hE0;
            16'd20151: data <= 8'h07;
            16'd20152: data <= 8'hE0;
            16'd20153: data <= 8'h07;
            16'd20154: data <= 8'hE0;
            16'd20155: data <= 8'h07;
            16'd20156: data <= 8'hE0;
            16'd20157: data <= 8'h07;
            16'd20158: data <= 8'hE0;
            16'd20159: data <= 8'h07;
            16'd20160: data <= 8'hFF;
            16'd20161: data <= 8'hFF;
            16'd20162: data <= 8'hE0;
            16'd20163: data <= 8'h07;
            16'd20164: data <= 8'hE0;
            16'd20165: data <= 8'h07;
            16'd20166: data <= 8'hE0;
            16'd20167: data <= 8'h07;
            16'd20168: data <= 8'hE0;
            16'd20169: data <= 8'h07;
            16'd20170: data <= 8'hE0;
            16'd20171: data <= 8'h07;
            16'd20172: data <= 8'hE0;
            16'd20173: data <= 8'h07;
            16'd20174: data <= 8'hE0;
            16'd20175: data <= 8'h07;
            16'd20176: data <= 8'hE0;
            16'd20177: data <= 8'h07;
            16'd20178: data <= 8'hE0;
            16'd20179: data <= 8'h07;
            16'd20180: data <= 8'hE0;
            16'd20181: data <= 8'h07;
            16'd20182: data <= 8'hE0;
            16'd20183: data <= 8'h07;
            16'd20184: data <= 8'hE0;
            16'd20185: data <= 8'h07;
            16'd20186: data <= 8'hE0;
            16'd20187: data <= 8'h07;
            16'd20188: data <= 8'hE0;
            16'd20189: data <= 8'h07;
            16'd20190: data <= 8'hE0;
            16'd20191: data <= 8'h07;
            16'd20192: data <= 8'hE0;
            16'd20193: data <= 8'h07;
            16'd20194: data <= 8'hE0;
            16'd20195: data <= 8'h07;
            16'd20196: data <= 8'hE0;
            16'd20197: data <= 8'h07;
            16'd20198: data <= 8'hE0;
            16'd20199: data <= 8'h07;
            16'd20200: data <= 8'hFF;
            16'd20201: data <= 8'hFF;
            16'd20202: data <= 8'hE0;
            16'd20203: data <= 8'h07;
            16'd20204: data <= 8'hE0;
            16'd20205: data <= 8'h07;
            16'd20206: data <= 8'hE0;
            16'd20207: data <= 8'h07;
            16'd20208: data <= 8'hE0;
            16'd20209: data <= 8'h07;
            16'd20210: data <= 8'hE0;
            16'd20211: data <= 8'h07;
            16'd20212: data <= 8'hE0;
            16'd20213: data <= 8'h07;
            16'd20214: data <= 8'hE0;
            16'd20215: data <= 8'h07;
            16'd20216: data <= 8'hE0;
            16'd20217: data <= 8'h07;
            16'd20218: data <= 8'hE0;
            16'd20219: data <= 8'h07;
            16'd20220: data <= 8'hE0;
            16'd20221: data <= 8'h07;
            16'd20222: data <= 8'hE0;
            16'd20223: data <= 8'h07;
            16'd20224: data <= 8'hE0;
            16'd20225: data <= 8'h07;
            16'd20226: data <= 8'hE0;
            16'd20227: data <= 8'h07;
            16'd20228: data <= 8'hE0;
            16'd20229: data <= 8'h07;
            16'd20230: data <= 8'hE0;
            16'd20231: data <= 8'h07;
            16'd20232: data <= 8'hE0;
            16'd20233: data <= 8'h07;
            16'd20234: data <= 8'hE0;
            16'd20235: data <= 8'h07;
            16'd20236: data <= 8'hE0;
            16'd20237: data <= 8'h07;
            16'd20238: data <= 8'hE0;
            16'd20239: data <= 8'h07;
            16'd20240: data <= 8'hFF;
            16'd20241: data <= 8'hFF;
            16'd20242: data <= 8'hE0;
            16'd20243: data <= 8'h07;
            16'd20244: data <= 8'hE0;
            16'd20245: data <= 8'h07;
            16'd20246: data <= 8'hE0;
            16'd20247: data <= 8'h07;
            16'd20248: data <= 8'hE0;
            16'd20249: data <= 8'h07;
            16'd20250: data <= 8'hE0;
            16'd20251: data <= 8'h07;
            16'd20252: data <= 8'hE0;
            16'd20253: data <= 8'h07;
            16'd20254: data <= 8'hE0;
            16'd20255: data <= 8'h07;
            16'd20256: data <= 8'hE0;
            16'd20257: data <= 8'h07;
            16'd20258: data <= 8'hE0;
            16'd20259: data <= 8'h07;
            16'd20260: data <= 8'hE0;
            16'd20261: data <= 8'h07;
            16'd20262: data <= 8'hE0;
            16'd20263: data <= 8'h07;
            16'd20264: data <= 8'hE0;
            16'd20265: data <= 8'h07;
            16'd20266: data <= 8'hE0;
            16'd20267: data <= 8'h07;
            16'd20268: data <= 8'hE0;
            16'd20269: data <= 8'h07;
            16'd20270: data <= 8'hE0;
            16'd20271: data <= 8'h07;
            16'd20272: data <= 8'hE0;
            16'd20273: data <= 8'h07;
            16'd20274: data <= 8'hE0;
            16'd20275: data <= 8'h07;
            16'd20276: data <= 8'hE0;
            16'd20277: data <= 8'h07;
            16'd20278: data <= 8'hE0;
            16'd20279: data <= 8'h07;
            16'd20280: data <= 8'hFF;
            16'd20281: data <= 8'hFF;
            16'd20282: data <= 8'hE0;
            16'd20283: data <= 8'h07;
            16'd20284: data <= 8'hE0;
            16'd20285: data <= 8'h07;
            16'd20286: data <= 8'hE0;
            16'd20287: data <= 8'h07;
            16'd20288: data <= 8'hE0;
            16'd20289: data <= 8'h07;
            16'd20290: data <= 8'hE0;
            16'd20291: data <= 8'h07;
            16'd20292: data <= 8'hE0;
            16'd20293: data <= 8'h07;
            16'd20294: data <= 8'hE0;
            16'd20295: data <= 8'h07;
            16'd20296: data <= 8'hE0;
            16'd20297: data <= 8'h07;
            16'd20298: data <= 8'hE0;
            16'd20299: data <= 8'h07;
            16'd20300: data <= 8'hE0;
            16'd20301: data <= 8'h07;
            16'd20302: data <= 8'hE0;
            16'd20303: data <= 8'h07;
            16'd20304: data <= 8'hE0;
            16'd20305: data <= 8'h07;
            16'd20306: data <= 8'hE0;
            16'd20307: data <= 8'h07;
            16'd20308: data <= 8'hE0;
            16'd20309: data <= 8'h07;
            16'd20310: data <= 8'hE0;
            16'd20311: data <= 8'h07;
            16'd20312: data <= 8'hE0;
            16'd20313: data <= 8'h07;
            16'd20314: data <= 8'hE0;
            16'd20315: data <= 8'h07;
            16'd20316: data <= 8'hE0;
            16'd20317: data <= 8'h07;
            16'd20318: data <= 8'hE0;
            16'd20319: data <= 8'h07;
            16'd20320: data <= 8'hFF;
            16'd20321: data <= 8'hFF;
            16'd20322: data <= 8'hE0;
            16'd20323: data <= 8'h07;
            16'd20324: data <= 8'hE0;
            16'd20325: data <= 8'h07;
            16'd20326: data <= 8'hE0;
            16'd20327: data <= 8'h07;
            16'd20328: data <= 8'hE0;
            16'd20329: data <= 8'h07;
            16'd20330: data <= 8'hE0;
            16'd20331: data <= 8'h07;
            16'd20332: data <= 8'hE0;
            16'd20333: data <= 8'h07;
            16'd20334: data <= 8'hE0;
            16'd20335: data <= 8'h07;
            16'd20336: data <= 8'hE0;
            16'd20337: data <= 8'h07;
            16'd20338: data <= 8'hE0;
            16'd20339: data <= 8'h07;
            16'd20340: data <= 8'hE0;
            16'd20341: data <= 8'h07;
            16'd20342: data <= 8'hE0;
            16'd20343: data <= 8'h07;
            16'd20344: data <= 8'hE0;
            16'd20345: data <= 8'h07;
            16'd20346: data <= 8'hE0;
            16'd20347: data <= 8'h07;
            16'd20348: data <= 8'hE0;
            16'd20349: data <= 8'h07;
            16'd20350: data <= 8'hE0;
            16'd20351: data <= 8'h07;
            16'd20352: data <= 8'hE0;
            16'd20353: data <= 8'h07;
            16'd20354: data <= 8'hE0;
            16'd20355: data <= 8'h07;
            16'd20356: data <= 8'hE0;
            16'd20357: data <= 8'h07;
            16'd20358: data <= 8'hE0;
            16'd20359: data <= 8'h07;
            16'd20360: data <= 8'hFF;
            16'd20361: data <= 8'hFF;
            16'd20362: data <= 8'hE0;
            16'd20363: data <= 8'h07;
            16'd20364: data <= 8'hE0;
            16'd20365: data <= 8'h07;
            16'd20366: data <= 8'hE0;
            16'd20367: data <= 8'h07;
            16'd20368: data <= 8'hE0;
            16'd20369: data <= 8'h07;
            16'd20370: data <= 8'hE0;
            16'd20371: data <= 8'h07;
            16'd20372: data <= 8'hE0;
            16'd20373: data <= 8'h07;
            16'd20374: data <= 8'hE0;
            16'd20375: data <= 8'h07;
            16'd20376: data <= 8'hE0;
            16'd20377: data <= 8'h07;
            16'd20378: data <= 8'hE0;
            16'd20379: data <= 8'h07;
            16'd20380: data <= 8'hE0;
            16'd20381: data <= 8'h07;
            16'd20382: data <= 8'hE0;
            16'd20383: data <= 8'h07;
            16'd20384: data <= 8'hE0;
            16'd20385: data <= 8'h07;
            16'd20386: data <= 8'hE0;
            16'd20387: data <= 8'h07;
            16'd20388: data <= 8'hE0;
            16'd20389: data <= 8'h07;
            16'd20390: data <= 8'hE0;
            16'd20391: data <= 8'h07;
            16'd20392: data <= 8'hE0;
            16'd20393: data <= 8'h07;
            16'd20394: data <= 8'hE0;
            16'd20395: data <= 8'h07;
            16'd20396: data <= 8'hE0;
            16'd20397: data <= 8'h07;
            16'd20398: data <= 8'hE0;
            16'd20399: data <= 8'h07;
            16'd20400: data <= 8'hFF;
            16'd20401: data <= 8'hFF;
            16'd20402: data <= 8'hE0;
            16'd20403: data <= 8'h07;
            16'd20404: data <= 8'hE0;
            16'd20405: data <= 8'h07;
            16'd20406: data <= 8'hE0;
            16'd20407: data <= 8'h07;
            16'd20408: data <= 8'hE0;
            16'd20409: data <= 8'h07;
            16'd20410: data <= 8'hE0;
            16'd20411: data <= 8'h07;
            16'd20412: data <= 8'hE0;
            16'd20413: data <= 8'h07;
            16'd20414: data <= 8'hE0;
            16'd20415: data <= 8'h07;
            16'd20416: data <= 8'hE0;
            16'd20417: data <= 8'h07;
            16'd20418: data <= 8'hE0;
            16'd20419: data <= 8'h07;
            16'd20420: data <= 8'hE0;
            16'd20421: data <= 8'h07;
            16'd20422: data <= 8'hE0;
            16'd20423: data <= 8'h07;
            16'd20424: data <= 8'hE0;
            16'd20425: data <= 8'h07;
            16'd20426: data <= 8'hE0;
            16'd20427: data <= 8'h07;
            16'd20428: data <= 8'hE0;
            16'd20429: data <= 8'h07;
            16'd20430: data <= 8'hE0;
            16'd20431: data <= 8'h07;
            16'd20432: data <= 8'hE0;
            16'd20433: data <= 8'h07;
            16'd20434: data <= 8'hE0;
            16'd20435: data <= 8'h07;
            16'd20436: data <= 8'hE0;
            16'd20437: data <= 8'h07;
            16'd20438: data <= 8'hE0;
            16'd20439: data <= 8'h07;
            16'd20440: data <= 8'hFF;
            16'd20441: data <= 8'hFF;
            16'd20442: data <= 8'hE0;
            16'd20443: data <= 8'h07;
            16'd20444: data <= 8'hE0;
            16'd20445: data <= 8'h07;
            16'd20446: data <= 8'hE0;
            16'd20447: data <= 8'h07;
            16'd20448: data <= 8'hE0;
            16'd20449: data <= 8'h07;
            16'd20450: data <= 8'hE0;
            16'd20451: data <= 8'h07;
            16'd20452: data <= 8'hE0;
            16'd20453: data <= 8'h07;
            16'd20454: data <= 8'hE0;
            16'd20455: data <= 8'h07;
            16'd20456: data <= 8'hE0;
            16'd20457: data <= 8'h07;
            16'd20458: data <= 8'hE0;
            16'd20459: data <= 8'h07;
            16'd20460: data <= 8'hE0;
            16'd20461: data <= 8'h07;
            16'd20462: data <= 8'hE0;
            16'd20463: data <= 8'h07;
            16'd20464: data <= 8'hE0;
            16'd20465: data <= 8'h07;
            16'd20466: data <= 8'hE0;
            16'd20467: data <= 8'h07;
            16'd20468: data <= 8'hE0;
            16'd20469: data <= 8'h07;
            16'd20470: data <= 8'hE0;
            16'd20471: data <= 8'h07;
            16'd20472: data <= 8'hE0;
            16'd20473: data <= 8'h07;
            16'd20474: data <= 8'hE0;
            16'd20475: data <= 8'h07;
            16'd20476: data <= 8'hE0;
            16'd20477: data <= 8'h07;
            16'd20478: data <= 8'hE0;
            16'd20479: data <= 8'h07;
            16'd20480: data <= 8'hFF;
            16'd20481: data <= 8'hFF;
            16'd20482: data <= 8'hE0;
            16'd20483: data <= 8'h07;
            16'd20484: data <= 8'hE0;
            16'd20485: data <= 8'h07;
            16'd20486: data <= 8'hE0;
            16'd20487: data <= 8'h07;
            16'd20488: data <= 8'hE0;
            16'd20489: data <= 8'h07;
            16'd20490: data <= 8'hE0;
            16'd20491: data <= 8'h07;
            16'd20492: data <= 8'hE0;
            16'd20493: data <= 8'h07;
            16'd20494: data <= 8'hE0;
            16'd20495: data <= 8'h07;
            16'd20496: data <= 8'hE0;
            16'd20497: data <= 8'h07;
            16'd20498: data <= 8'hE0;
            16'd20499: data <= 8'h07;
            16'd20500: data <= 8'hE0;
            16'd20501: data <= 8'h07;
            16'd20502: data <= 8'hE0;
            16'd20503: data <= 8'h07;
            16'd20504: data <= 8'hE0;
            16'd20505: data <= 8'h07;
            16'd20506: data <= 8'hE0;
            16'd20507: data <= 8'h07;
            16'd20508: data <= 8'hE0;
            16'd20509: data <= 8'h07;
            16'd20510: data <= 8'hE0;
            16'd20511: data <= 8'h07;
            16'd20512: data <= 8'hE0;
            16'd20513: data <= 8'h07;
            16'd20514: data <= 8'hE0;
            16'd20515: data <= 8'h07;
            16'd20516: data <= 8'hE0;
            16'd20517: data <= 8'h07;
            16'd20518: data <= 8'hE0;
            16'd20519: data <= 8'h07;
            16'd20520: data <= 8'hFF;
            16'd20521: data <= 8'hFF;
            16'd20522: data <= 8'hE0;
            16'd20523: data <= 8'h07;
            16'd20524: data <= 8'hE0;
            16'd20525: data <= 8'h07;
            16'd20526: data <= 8'hE0;
            16'd20527: data <= 8'h07;
            16'd20528: data <= 8'hE0;
            16'd20529: data <= 8'h07;
            16'd20530: data <= 8'hE0;
            16'd20531: data <= 8'h07;
            16'd20532: data <= 8'hE0;
            16'd20533: data <= 8'h07;
            16'd20534: data <= 8'hE0;
            16'd20535: data <= 8'h07;
            16'd20536: data <= 8'hE0;
            16'd20537: data <= 8'h07;
            16'd20538: data <= 8'hE0;
            16'd20539: data <= 8'h07;
            16'd20540: data <= 8'hE0;
            16'd20541: data <= 8'h07;
            16'd20542: data <= 8'hE0;
            16'd20543: data <= 8'h07;
            16'd20544: data <= 8'hE0;
            16'd20545: data <= 8'h07;
            16'd20546: data <= 8'hE0;
            16'd20547: data <= 8'h07;
            16'd20548: data <= 8'hE0;
            16'd20549: data <= 8'h07;
            16'd20550: data <= 8'hE0;
            16'd20551: data <= 8'h07;
            16'd20552: data <= 8'hE0;
            16'd20553: data <= 8'h07;
            16'd20554: data <= 8'hE0;
            16'd20555: data <= 8'h07;
            16'd20556: data <= 8'hE0;
            16'd20557: data <= 8'h07;
            16'd20558: data <= 8'hE0;
            16'd20559: data <= 8'h07;
            16'd20560: data <= 8'hFF;
            16'd20561: data <= 8'hFF;
            16'd20562: data <= 8'hE0;
            16'd20563: data <= 8'h07;
            16'd20564: data <= 8'hE0;
            16'd20565: data <= 8'h07;
            16'd20566: data <= 8'hE0;
            16'd20567: data <= 8'h07;
            16'd20568: data <= 8'hE0;
            16'd20569: data <= 8'h07;
            16'd20570: data <= 8'hE0;
            16'd20571: data <= 8'h07;
            16'd20572: data <= 8'hE0;
            16'd20573: data <= 8'h07;
            16'd20574: data <= 8'hE0;
            16'd20575: data <= 8'h07;
            16'd20576: data <= 8'hE0;
            16'd20577: data <= 8'h07;
            16'd20578: data <= 8'hE0;
            16'd20579: data <= 8'h07;
            16'd20580: data <= 8'hE0;
            16'd20581: data <= 8'h07;
            16'd20582: data <= 8'hE0;
            16'd20583: data <= 8'h07;
            16'd20584: data <= 8'hE0;
            16'd20585: data <= 8'h07;
            16'd20586: data <= 8'hE0;
            16'd20587: data <= 8'h07;
            16'd20588: data <= 8'hE0;
            16'd20589: data <= 8'h07;
            16'd20590: data <= 8'hE0;
            16'd20591: data <= 8'h07;
            16'd20592: data <= 8'hE0;
            16'd20593: data <= 8'h07;
            16'd20594: data <= 8'hE0;
            16'd20595: data <= 8'h07;
            16'd20596: data <= 8'hE0;
            16'd20597: data <= 8'h07;
            16'd20598: data <= 8'hE0;
            16'd20599: data <= 8'h07;
            16'd20600: data <= 8'hFF;
            16'd20601: data <= 8'hFF;
            16'd20602: data <= 8'hE0;
            16'd20603: data <= 8'h07;
            16'd20604: data <= 8'hE0;
            16'd20605: data <= 8'h07;
            16'd20606: data <= 8'hE0;
            16'd20607: data <= 8'h07;
            16'd20608: data <= 8'hE0;
            16'd20609: data <= 8'h07;
            16'd20610: data <= 8'hE0;
            16'd20611: data <= 8'h07;
            16'd20612: data <= 8'hE0;
            16'd20613: data <= 8'h07;
            16'd20614: data <= 8'hE0;
            16'd20615: data <= 8'h07;
            16'd20616: data <= 8'hE0;
            16'd20617: data <= 8'h07;
            16'd20618: data <= 8'hE0;
            16'd20619: data <= 8'h07;
            16'd20620: data <= 8'hE0;
            16'd20621: data <= 8'h07;
            16'd20622: data <= 8'hE0;
            16'd20623: data <= 8'h07;
            16'd20624: data <= 8'hE0;
            16'd20625: data <= 8'h07;
            16'd20626: data <= 8'hE0;
            16'd20627: data <= 8'h07;
            16'd20628: data <= 8'hE0;
            16'd20629: data <= 8'h07;
            16'd20630: data <= 8'hE0;
            16'd20631: data <= 8'h07;
            16'd20632: data <= 8'hE0;
            16'd20633: data <= 8'h07;
            16'd20634: data <= 8'hE0;
            16'd20635: data <= 8'h07;
            16'd20636: data <= 8'hE0;
            16'd20637: data <= 8'h07;
            16'd20638: data <= 8'hE0;
            16'd20639: data <= 8'h07;
            16'd20640: data <= 8'hFF;
            16'd20641: data <= 8'hFF;
            16'd20642: data <= 8'hE0;
            16'd20643: data <= 8'h07;
            16'd20644: data <= 8'hE0;
            16'd20645: data <= 8'h07;
            16'd20646: data <= 8'hE0;
            16'd20647: data <= 8'h07;
            16'd20648: data <= 8'hE0;
            16'd20649: data <= 8'h07;
            16'd20650: data <= 8'hE0;
            16'd20651: data <= 8'h07;
            16'd20652: data <= 8'hE0;
            16'd20653: data <= 8'h07;
            16'd20654: data <= 8'hE0;
            16'd20655: data <= 8'h07;
            16'd20656: data <= 8'hE0;
            16'd20657: data <= 8'h07;
            16'd20658: data <= 8'hE0;
            16'd20659: data <= 8'h07;
            16'd20660: data <= 8'hE0;
            16'd20661: data <= 8'h07;
            16'd20662: data <= 8'hE0;
            16'd20663: data <= 8'h07;
            16'd20664: data <= 8'hE0;
            16'd20665: data <= 8'h07;
            16'd20666: data <= 8'hE0;
            16'd20667: data <= 8'h07;
            16'd20668: data <= 8'hE0;
            16'd20669: data <= 8'h07;
            16'd20670: data <= 8'hE0;
            16'd20671: data <= 8'h07;
            16'd20672: data <= 8'hE0;
            16'd20673: data <= 8'h07;
            16'd20674: data <= 8'hE0;
            16'd20675: data <= 8'h07;
            16'd20676: data <= 8'hE0;
            16'd20677: data <= 8'h07;
            16'd20678: data <= 8'hE0;
            16'd20679: data <= 8'h07;
            16'd20680: data <= 8'hFF;
            16'd20681: data <= 8'hFF;
            16'd20682: data <= 8'hE0;
            16'd20683: data <= 8'h07;
            16'd20684: data <= 8'hE0;
            16'd20685: data <= 8'h07;
            16'd20686: data <= 8'hE0;
            16'd20687: data <= 8'h07;
            16'd20688: data <= 8'hE0;
            16'd20689: data <= 8'h07;
            16'd20690: data <= 8'hE0;
            16'd20691: data <= 8'h07;
            16'd20692: data <= 8'hE0;
            16'd20693: data <= 8'h07;
            16'd20694: data <= 8'hE0;
            16'd20695: data <= 8'h07;
            16'd20696: data <= 8'hE0;
            16'd20697: data <= 8'h07;
            16'd20698: data <= 8'hE0;
            16'd20699: data <= 8'h07;
            16'd20700: data <= 8'hE0;
            16'd20701: data <= 8'h07;
            16'd20702: data <= 8'hE0;
            16'd20703: data <= 8'h07;
            16'd20704: data <= 8'hE0;
            16'd20705: data <= 8'h07;
            16'd20706: data <= 8'hE0;
            16'd20707: data <= 8'h07;
            16'd20708: data <= 8'hE0;
            16'd20709: data <= 8'h07;
            16'd20710: data <= 8'hE0;
            16'd20711: data <= 8'h07;
            16'd20712: data <= 8'hE0;
            16'd20713: data <= 8'h07;
            16'd20714: data <= 8'hE0;
            16'd20715: data <= 8'h07;
            16'd20716: data <= 8'hE0;
            16'd20717: data <= 8'h07;
            16'd20718: data <= 8'hE0;
            16'd20719: data <= 8'h07;
            16'd20720: data <= 8'hFF;
            16'd20721: data <= 8'hFF;
            16'd20722: data <= 8'hE0;
            16'd20723: data <= 8'h07;
            16'd20724: data <= 8'hE0;
            16'd20725: data <= 8'h07;
            16'd20726: data <= 8'hE0;
            16'd20727: data <= 8'h07;
            16'd20728: data <= 8'hE0;
            16'd20729: data <= 8'h07;
            16'd20730: data <= 8'hE0;
            16'd20731: data <= 8'h07;
            16'd20732: data <= 8'hE0;
            16'd20733: data <= 8'h07;
            16'd20734: data <= 8'hE0;
            16'd20735: data <= 8'h07;
            16'd20736: data <= 8'hE0;
            16'd20737: data <= 8'h07;
            16'd20738: data <= 8'hE0;
            16'd20739: data <= 8'h07;
            16'd20740: data <= 8'hE0;
            16'd20741: data <= 8'h07;
            16'd20742: data <= 8'hE0;
            16'd20743: data <= 8'h07;
            16'd20744: data <= 8'hE0;
            16'd20745: data <= 8'h07;
            16'd20746: data <= 8'hE0;
            16'd20747: data <= 8'h07;
            16'd20748: data <= 8'hE0;
            16'd20749: data <= 8'h07;
            16'd20750: data <= 8'hE0;
            16'd20751: data <= 8'h07;
            16'd20752: data <= 8'hE0;
            16'd20753: data <= 8'h07;
            16'd20754: data <= 8'hE0;
            16'd20755: data <= 8'h07;
            16'd20756: data <= 8'hE0;
            16'd20757: data <= 8'h07;
            16'd20758: data <= 8'hE0;
            16'd20759: data <= 8'h07;
            16'd20760: data <= 8'hFF;
            16'd20761: data <= 8'hFF;
            16'd20762: data <= 8'hE0;
            16'd20763: data <= 8'h07;
            16'd20764: data <= 8'hE0;
            16'd20765: data <= 8'h07;
            16'd20766: data <= 8'hE0;
            16'd20767: data <= 8'h07;
            16'd20768: data <= 8'hE0;
            16'd20769: data <= 8'h07;
            16'd20770: data <= 8'hE0;
            16'd20771: data <= 8'h07;
            16'd20772: data <= 8'hE0;
            16'd20773: data <= 8'h07;
            16'd20774: data <= 8'hE0;
            16'd20775: data <= 8'h07;
            16'd20776: data <= 8'hE0;
            16'd20777: data <= 8'h07;
            16'd20778: data <= 8'hE0;
            16'd20779: data <= 8'h07;
            16'd20780: data <= 8'hE0;
            16'd20781: data <= 8'h07;
            16'd20782: data <= 8'hE0;
            16'd20783: data <= 8'h07;
            16'd20784: data <= 8'hE0;
            16'd20785: data <= 8'h07;
            16'd20786: data <= 8'hE0;
            16'd20787: data <= 8'h07;
            16'd20788: data <= 8'hE0;
            16'd20789: data <= 8'h07;
            16'd20790: data <= 8'hE0;
            16'd20791: data <= 8'h07;
            16'd20792: data <= 8'hE0;
            16'd20793: data <= 8'h07;
            16'd20794: data <= 8'hE0;
            16'd20795: data <= 8'h07;
            16'd20796: data <= 8'hE0;
            16'd20797: data <= 8'h07;
            16'd20798: data <= 8'hE0;
            16'd20799: data <= 8'h07;
            16'd20800: data <= 8'hFF;
            16'd20801: data <= 8'hFF;
            16'd20802: data <= 8'hE0;
            16'd20803: data <= 8'h07;
            16'd20804: data <= 8'hE0;
            16'd20805: data <= 8'h07;
            16'd20806: data <= 8'hE0;
            16'd20807: data <= 8'h07;
            16'd20808: data <= 8'hE0;
            16'd20809: data <= 8'h07;
            16'd20810: data <= 8'hE0;
            16'd20811: data <= 8'h07;
            16'd20812: data <= 8'hE0;
            16'd20813: data <= 8'h07;
            16'd20814: data <= 8'hE0;
            16'd20815: data <= 8'h07;
            16'd20816: data <= 8'hE0;
            16'd20817: data <= 8'h07;
            16'd20818: data <= 8'hE0;
            16'd20819: data <= 8'h07;
            16'd20820: data <= 8'hE0;
            16'd20821: data <= 8'h07;
            16'd20822: data <= 8'hE0;
            16'd20823: data <= 8'h07;
            16'd20824: data <= 8'hE0;
            16'd20825: data <= 8'h07;
            16'd20826: data <= 8'hE0;
            16'd20827: data <= 8'h07;
            16'd20828: data <= 8'hE0;
            16'd20829: data <= 8'h07;
            16'd20830: data <= 8'hE0;
            16'd20831: data <= 8'h07;
            16'd20832: data <= 8'hE0;
            16'd20833: data <= 8'h07;
            16'd20834: data <= 8'hE0;
            16'd20835: data <= 8'h07;
            16'd20836: data <= 8'hE0;
            16'd20837: data <= 8'h07;
            16'd20838: data <= 8'hE0;
            16'd20839: data <= 8'h07;
            16'd20840: data <= 8'hFF;
            16'd20841: data <= 8'hFF;
            16'd20842: data <= 8'hE0;
            16'd20843: data <= 8'h07;
            16'd20844: data <= 8'hE0;
            16'd20845: data <= 8'h07;
            16'd20846: data <= 8'hE0;
            16'd20847: data <= 8'h07;
            16'd20848: data <= 8'hE0;
            16'd20849: data <= 8'h07;
            16'd20850: data <= 8'hE0;
            16'd20851: data <= 8'h07;
            16'd20852: data <= 8'hE0;
            16'd20853: data <= 8'h07;
            16'd20854: data <= 8'hE0;
            16'd20855: data <= 8'h07;
            16'd20856: data <= 8'hE0;
            16'd20857: data <= 8'h07;
            16'd20858: data <= 8'hE0;
            16'd20859: data <= 8'h07;
            16'd20860: data <= 8'hE0;
            16'd20861: data <= 8'h07;
            16'd20862: data <= 8'hE0;
            16'd20863: data <= 8'h07;
            16'd20864: data <= 8'hE0;
            16'd20865: data <= 8'h07;
            16'd20866: data <= 8'hE0;
            16'd20867: data <= 8'h07;
            16'd20868: data <= 8'hE0;
            16'd20869: data <= 8'h07;
            16'd20870: data <= 8'hE0;
            16'd20871: data <= 8'h07;
            16'd20872: data <= 8'hE0;
            16'd20873: data <= 8'h07;
            16'd20874: data <= 8'hE0;
            16'd20875: data <= 8'h07;
            16'd20876: data <= 8'hE0;
            16'd20877: data <= 8'h07;
            16'd20878: data <= 8'hE0;
            16'd20879: data <= 8'h07;
            16'd20880: data <= 8'hFF;
            16'd20881: data <= 8'hFF;
            16'd20882: data <= 8'hE0;
            16'd20883: data <= 8'h07;
            16'd20884: data <= 8'hE0;
            16'd20885: data <= 8'h07;
            16'd20886: data <= 8'hE0;
            16'd20887: data <= 8'h07;
            16'd20888: data <= 8'hE0;
            16'd20889: data <= 8'h07;
            16'd20890: data <= 8'hE0;
            16'd20891: data <= 8'h07;
            16'd20892: data <= 8'hE0;
            16'd20893: data <= 8'h07;
            16'd20894: data <= 8'hE0;
            16'd20895: data <= 8'h07;
            16'd20896: data <= 8'hE0;
            16'd20897: data <= 8'h07;
            16'd20898: data <= 8'hE0;
            16'd20899: data <= 8'h07;
            16'd20900: data <= 8'hE0;
            16'd20901: data <= 8'h07;
            16'd20902: data <= 8'hE0;
            16'd20903: data <= 8'h07;
            16'd20904: data <= 8'hE0;
            16'd20905: data <= 8'h07;
            16'd20906: data <= 8'hE0;
            16'd20907: data <= 8'h07;
            16'd20908: data <= 8'hE0;
            16'd20909: data <= 8'h07;
            16'd20910: data <= 8'hE0;
            16'd20911: data <= 8'h07;
            16'd20912: data <= 8'hE0;
            16'd20913: data <= 8'h07;
            16'd20914: data <= 8'hE0;
            16'd20915: data <= 8'h07;
            16'd20916: data <= 8'hE0;
            16'd20917: data <= 8'h07;
            16'd20918: data <= 8'hE0;
            16'd20919: data <= 8'h07;
            16'd20920: data <= 8'hFF;
            16'd20921: data <= 8'hFF;
            16'd20922: data <= 8'hE0;
            16'd20923: data <= 8'h07;
            16'd20924: data <= 8'hE0;
            16'd20925: data <= 8'h07;
            16'd20926: data <= 8'hE0;
            16'd20927: data <= 8'h07;
            16'd20928: data <= 8'hE0;
            16'd20929: data <= 8'h07;
            16'd20930: data <= 8'hE0;
            16'd20931: data <= 8'h07;
            16'd20932: data <= 8'hE0;
            16'd20933: data <= 8'h07;
            16'd20934: data <= 8'hE0;
            16'd20935: data <= 8'h07;
            16'd20936: data <= 8'hE0;
            16'd20937: data <= 8'h07;
            16'd20938: data <= 8'hE0;
            16'd20939: data <= 8'h07;
            16'd20940: data <= 8'hE0;
            16'd20941: data <= 8'h07;
            16'd20942: data <= 8'hE0;
            16'd20943: data <= 8'h07;
            16'd20944: data <= 8'hE0;
            16'd20945: data <= 8'h07;
            16'd20946: data <= 8'hE0;
            16'd20947: data <= 8'h07;
            16'd20948: data <= 8'hE0;
            16'd20949: data <= 8'h07;
            16'd20950: data <= 8'hE0;
            16'd20951: data <= 8'h07;
            16'd20952: data <= 8'hE0;
            16'd20953: data <= 8'h07;
            16'd20954: data <= 8'hE0;
            16'd20955: data <= 8'h07;
            16'd20956: data <= 8'hE0;
            16'd20957: data <= 8'h07;
            16'd20958: data <= 8'hE0;
            16'd20959: data <= 8'h07;
            16'd20960: data <= 8'hFF;
            16'd20961: data <= 8'hFF;
            16'd20962: data <= 8'hE0;
            16'd20963: data <= 8'h07;
            16'd20964: data <= 8'hE0;
            16'd20965: data <= 8'h07;
            16'd20966: data <= 8'hE0;
            16'd20967: data <= 8'h07;
            16'd20968: data <= 8'hE0;
            16'd20969: data <= 8'h07;
            16'd20970: data <= 8'hE0;
            16'd20971: data <= 8'h07;
            16'd20972: data <= 8'hE0;
            16'd20973: data <= 8'h07;
            16'd20974: data <= 8'hE0;
            16'd20975: data <= 8'h07;
            16'd20976: data <= 8'hE0;
            16'd20977: data <= 8'h07;
            16'd20978: data <= 8'hE0;
            16'd20979: data <= 8'h07;
            16'd20980: data <= 8'hE0;
            16'd20981: data <= 8'h07;
            16'd20982: data <= 8'hE0;
            16'd20983: data <= 8'h07;
            16'd20984: data <= 8'hE0;
            16'd20985: data <= 8'h07;
            16'd20986: data <= 8'hE0;
            16'd20987: data <= 8'h07;
            16'd20988: data <= 8'hE0;
            16'd20989: data <= 8'h07;
            16'd20990: data <= 8'hE0;
            16'd20991: data <= 8'h07;
            16'd20992: data <= 8'hE0;
            16'd20993: data <= 8'h07;
            16'd20994: data <= 8'hE0;
            16'd20995: data <= 8'h07;
            16'd20996: data <= 8'hE0;
            16'd20997: data <= 8'h07;
            16'd20998: data <= 8'hE0;
            16'd20999: data <= 8'h07;
            16'd21000: data <= 8'hFF;
            16'd21001: data <= 8'hFF;
            16'd21002: data <= 8'hE0;
            16'd21003: data <= 8'h07;
            16'd21004: data <= 8'hE0;
            16'd21005: data <= 8'h07;
            16'd21006: data <= 8'hE0;
            16'd21007: data <= 8'h07;
            16'd21008: data <= 8'hE0;
            16'd21009: data <= 8'h07;
            16'd21010: data <= 8'hE0;
            16'd21011: data <= 8'h07;
            16'd21012: data <= 8'hE0;
            16'd21013: data <= 8'h07;
            16'd21014: data <= 8'hE0;
            16'd21015: data <= 8'h07;
            16'd21016: data <= 8'hE0;
            16'd21017: data <= 8'h07;
            16'd21018: data <= 8'hE0;
            16'd21019: data <= 8'h07;
            16'd21020: data <= 8'hE0;
            16'd21021: data <= 8'h07;
            16'd21022: data <= 8'hE0;
            16'd21023: data <= 8'h07;
            16'd21024: data <= 8'hE0;
            16'd21025: data <= 8'h07;
            16'd21026: data <= 8'hE0;
            16'd21027: data <= 8'h07;
            16'd21028: data <= 8'hE0;
            16'd21029: data <= 8'h07;
            16'd21030: data <= 8'hE0;
            16'd21031: data <= 8'h07;
            16'd21032: data <= 8'hE0;
            16'd21033: data <= 8'h07;
            16'd21034: data <= 8'hE0;
            16'd21035: data <= 8'h07;
            16'd21036: data <= 8'hE0;
            16'd21037: data <= 8'h07;
            16'd21038: data <= 8'hE0;
            16'd21039: data <= 8'h07;
            16'd21040: data <= 8'hFF;
            16'd21041: data <= 8'hFF;
            16'd21042: data <= 8'hE0;
            16'd21043: data <= 8'h07;
            16'd21044: data <= 8'hE0;
            16'd21045: data <= 8'h07;
            16'd21046: data <= 8'hE0;
            16'd21047: data <= 8'h07;
            16'd21048: data <= 8'hE0;
            16'd21049: data <= 8'h07;
            16'd21050: data <= 8'hE0;
            16'd21051: data <= 8'h07;
            16'd21052: data <= 8'hE0;
            16'd21053: data <= 8'h07;
            16'd21054: data <= 8'hE0;
            16'd21055: data <= 8'h07;
            16'd21056: data <= 8'hE0;
            16'd21057: data <= 8'h07;
            16'd21058: data <= 8'hE0;
            16'd21059: data <= 8'h07;
            16'd21060: data <= 8'hE0;
            16'd21061: data <= 8'h07;
            16'd21062: data <= 8'hE0;
            16'd21063: data <= 8'h07;
            16'd21064: data <= 8'hE0;
            16'd21065: data <= 8'h07;
            16'd21066: data <= 8'hE0;
            16'd21067: data <= 8'h07;
            16'd21068: data <= 8'hE0;
            16'd21069: data <= 8'h07;
            16'd21070: data <= 8'hE0;
            16'd21071: data <= 8'h07;
            16'd21072: data <= 8'hE0;
            16'd21073: data <= 8'h07;
            16'd21074: data <= 8'hE0;
            16'd21075: data <= 8'h07;
            16'd21076: data <= 8'hE0;
            16'd21077: data <= 8'h07;
            16'd21078: data <= 8'hE0;
            16'd21079: data <= 8'h07;
            16'd21080: data <= 8'hFF;
            16'd21081: data <= 8'hFF;
            16'd21082: data <= 8'hE0;
            16'd21083: data <= 8'h07;
            16'd21084: data <= 8'hE0;
            16'd21085: data <= 8'h07;
            16'd21086: data <= 8'hE0;
            16'd21087: data <= 8'h07;
            16'd21088: data <= 8'hE0;
            16'd21089: data <= 8'h07;
            16'd21090: data <= 8'hE0;
            16'd21091: data <= 8'h07;
            16'd21092: data <= 8'hE0;
            16'd21093: data <= 8'h07;
            16'd21094: data <= 8'hE0;
            16'd21095: data <= 8'h07;
            16'd21096: data <= 8'hE0;
            16'd21097: data <= 8'h07;
            16'd21098: data <= 8'hE0;
            16'd21099: data <= 8'h07;
            16'd21100: data <= 8'hE0;
            16'd21101: data <= 8'h07;
            16'd21102: data <= 8'hE0;
            16'd21103: data <= 8'h07;
            16'd21104: data <= 8'hE0;
            16'd21105: data <= 8'h07;
            16'd21106: data <= 8'hE0;
            16'd21107: data <= 8'h07;
            16'd21108: data <= 8'hE0;
            16'd21109: data <= 8'h07;
            16'd21110: data <= 8'hE0;
            16'd21111: data <= 8'h07;
            16'd21112: data <= 8'hE0;
            16'd21113: data <= 8'h07;
            16'd21114: data <= 8'hE0;
            16'd21115: data <= 8'h07;
            16'd21116: data <= 8'hE0;
            16'd21117: data <= 8'h07;
            16'd21118: data <= 8'hE0;
            16'd21119: data <= 8'h07;
            16'd21120: data <= 8'hFF;
            16'd21121: data <= 8'hFF;
            16'd21122: data <= 8'hE0;
            16'd21123: data <= 8'h07;
            16'd21124: data <= 8'hE0;
            16'd21125: data <= 8'h07;
            16'd21126: data <= 8'hE0;
            16'd21127: data <= 8'h07;
            16'd21128: data <= 8'hE0;
            16'd21129: data <= 8'h07;
            16'd21130: data <= 8'hE0;
            16'd21131: data <= 8'h07;
            16'd21132: data <= 8'hE0;
            16'd21133: data <= 8'h07;
            16'd21134: data <= 8'hE0;
            16'd21135: data <= 8'h07;
            16'd21136: data <= 8'hE0;
            16'd21137: data <= 8'h07;
            16'd21138: data <= 8'hE0;
            16'd21139: data <= 8'h07;
            16'd21140: data <= 8'hE0;
            16'd21141: data <= 8'h07;
            16'd21142: data <= 8'hE0;
            16'd21143: data <= 8'h07;
            16'd21144: data <= 8'hE0;
            16'd21145: data <= 8'h07;
            16'd21146: data <= 8'hE0;
            16'd21147: data <= 8'h07;
            16'd21148: data <= 8'hE0;
            16'd21149: data <= 8'h07;
            16'd21150: data <= 8'hE0;
            16'd21151: data <= 8'h07;
            16'd21152: data <= 8'hE0;
            16'd21153: data <= 8'h07;
            16'd21154: data <= 8'hE0;
            16'd21155: data <= 8'h07;
            16'd21156: data <= 8'hE0;
            16'd21157: data <= 8'h07;
            16'd21158: data <= 8'hE0;
            16'd21159: data <= 8'h07;
            16'd21160: data <= 8'hFF;
            16'd21161: data <= 8'hFF;
            16'd21162: data <= 8'hE0;
            16'd21163: data <= 8'h07;
            16'd21164: data <= 8'hE0;
            16'd21165: data <= 8'h07;
            16'd21166: data <= 8'hE0;
            16'd21167: data <= 8'h07;
            16'd21168: data <= 8'hE0;
            16'd21169: data <= 8'h07;
            16'd21170: data <= 8'hE0;
            16'd21171: data <= 8'h07;
            16'd21172: data <= 8'hE0;
            16'd21173: data <= 8'h07;
            16'd21174: data <= 8'hE0;
            16'd21175: data <= 8'h07;
            16'd21176: data <= 8'hE0;
            16'd21177: data <= 8'h07;
            16'd21178: data <= 8'hE0;
            16'd21179: data <= 8'h07;
            16'd21180: data <= 8'hE0;
            16'd21181: data <= 8'h07;
            16'd21182: data <= 8'hE0;
            16'd21183: data <= 8'h07;
            16'd21184: data <= 8'hE0;
            16'd21185: data <= 8'h07;
            16'd21186: data <= 8'hE0;
            16'd21187: data <= 8'h07;
            16'd21188: data <= 8'hE0;
            16'd21189: data <= 8'h07;
            16'd21190: data <= 8'hE0;
            16'd21191: data <= 8'h07;
            16'd21192: data <= 8'hE0;
            16'd21193: data <= 8'h07;
            16'd21194: data <= 8'hE0;
            16'd21195: data <= 8'h07;
            16'd21196: data <= 8'hE0;
            16'd21197: data <= 8'h07;
            16'd21198: data <= 8'hE0;
            16'd21199: data <= 8'h07;
            16'd21200: data <= 8'hFF;
            16'd21201: data <= 8'hFF;
            16'd21202: data <= 8'hE0;
            16'd21203: data <= 8'h07;
            16'd21204: data <= 8'hE0;
            16'd21205: data <= 8'h07;
            16'd21206: data <= 8'hE0;
            16'd21207: data <= 8'h07;
            16'd21208: data <= 8'hE0;
            16'd21209: data <= 8'h07;
            16'd21210: data <= 8'hE0;
            16'd21211: data <= 8'h07;
            16'd21212: data <= 8'hE0;
            16'd21213: data <= 8'h07;
            16'd21214: data <= 8'hE0;
            16'd21215: data <= 8'h07;
            16'd21216: data <= 8'hE0;
            16'd21217: data <= 8'h07;
            16'd21218: data <= 8'hE0;
            16'd21219: data <= 8'h07;
            16'd21220: data <= 8'hE0;
            16'd21221: data <= 8'h07;
            16'd21222: data <= 8'hE0;
            16'd21223: data <= 8'h07;
            16'd21224: data <= 8'hE0;
            16'd21225: data <= 8'h07;
            16'd21226: data <= 8'hE0;
            16'd21227: data <= 8'h07;
            16'd21228: data <= 8'hE0;
            16'd21229: data <= 8'h07;
            16'd21230: data <= 8'hE0;
            16'd21231: data <= 8'h07;
            16'd21232: data <= 8'hE0;
            16'd21233: data <= 8'h07;
            16'd21234: data <= 8'hE0;
            16'd21235: data <= 8'h07;
            16'd21236: data <= 8'hE0;
            16'd21237: data <= 8'h07;
            16'd21238: data <= 8'hE0;
            16'd21239: data <= 8'h07;
            16'd21240: data <= 8'hFF;
            16'd21241: data <= 8'hFF;
            16'd21242: data <= 8'hE0;
            16'd21243: data <= 8'h07;
            16'd21244: data <= 8'hE0;
            16'd21245: data <= 8'h07;
            16'd21246: data <= 8'hE0;
            16'd21247: data <= 8'h07;
            16'd21248: data <= 8'hE0;
            16'd21249: data <= 8'h07;
            16'd21250: data <= 8'hE0;
            16'd21251: data <= 8'h07;
            16'd21252: data <= 8'hE0;
            16'd21253: data <= 8'h07;
            16'd21254: data <= 8'hE0;
            16'd21255: data <= 8'h07;
            16'd21256: data <= 8'hE0;
            16'd21257: data <= 8'h07;
            16'd21258: data <= 8'hE0;
            16'd21259: data <= 8'h07;
            16'd21260: data <= 8'hE0;
            16'd21261: data <= 8'h07;
            16'd21262: data <= 8'hE0;
            16'd21263: data <= 8'h07;
            16'd21264: data <= 8'hE0;
            16'd21265: data <= 8'h07;
            16'd21266: data <= 8'hE0;
            16'd21267: data <= 8'h07;
            16'd21268: data <= 8'hE0;
            16'd21269: data <= 8'h07;
            16'd21270: data <= 8'hE0;
            16'd21271: data <= 8'h07;
            16'd21272: data <= 8'hE0;
            16'd21273: data <= 8'h07;
            16'd21274: data <= 8'hE0;
            16'd21275: data <= 8'h07;
            16'd21276: data <= 8'hE0;
            16'd21277: data <= 8'h07;
            16'd21278: data <= 8'hE0;
            16'd21279: data <= 8'h07;
            16'd21280: data <= 8'hFF;
            16'd21281: data <= 8'hFF;
            16'd21282: data <= 8'hE0;
            16'd21283: data <= 8'h07;
            16'd21284: data <= 8'hE0;
            16'd21285: data <= 8'h07;
            16'd21286: data <= 8'hE0;
            16'd21287: data <= 8'h07;
            16'd21288: data <= 8'hE0;
            16'd21289: data <= 8'h07;
            16'd21290: data <= 8'hE0;
            16'd21291: data <= 8'h07;
            16'd21292: data <= 8'hE0;
            16'd21293: data <= 8'h07;
            16'd21294: data <= 8'hE0;
            16'd21295: data <= 8'h07;
            16'd21296: data <= 8'hE0;
            16'd21297: data <= 8'h07;
            16'd21298: data <= 8'hE0;
            16'd21299: data <= 8'h07;
            16'd21300: data <= 8'hE0;
            16'd21301: data <= 8'h07;
            16'd21302: data <= 8'hE0;
            16'd21303: data <= 8'h07;
            16'd21304: data <= 8'hE0;
            16'd21305: data <= 8'h07;
            16'd21306: data <= 8'hE0;
            16'd21307: data <= 8'h07;
            16'd21308: data <= 8'hE0;
            16'd21309: data <= 8'h07;
            16'd21310: data <= 8'hE0;
            16'd21311: data <= 8'h07;
            16'd21312: data <= 8'hE0;
            16'd21313: data <= 8'h07;
            16'd21314: data <= 8'hE0;
            16'd21315: data <= 8'h07;
            16'd21316: data <= 8'hE0;
            16'd21317: data <= 8'h07;
            16'd21318: data <= 8'hE0;
            16'd21319: data <= 8'h07;
            16'd21320: data <= 8'hFF;
            16'd21321: data <= 8'hFF;
            16'd21322: data <= 8'hE0;
            16'd21323: data <= 8'h07;
            16'd21324: data <= 8'hE0;
            16'd21325: data <= 8'h07;
            16'd21326: data <= 8'hE0;
            16'd21327: data <= 8'h07;
            16'd21328: data <= 8'hE0;
            16'd21329: data <= 8'h07;
            16'd21330: data <= 8'hE0;
            16'd21331: data <= 8'h07;
            16'd21332: data <= 8'hE0;
            16'd21333: data <= 8'h07;
            16'd21334: data <= 8'hE0;
            16'd21335: data <= 8'h07;
            16'd21336: data <= 8'hE0;
            16'd21337: data <= 8'h07;
            16'd21338: data <= 8'hE0;
            16'd21339: data <= 8'h07;
            16'd21340: data <= 8'hE0;
            16'd21341: data <= 8'h07;
            16'd21342: data <= 8'hE0;
            16'd21343: data <= 8'h07;
            16'd21344: data <= 8'hE0;
            16'd21345: data <= 8'h07;
            16'd21346: data <= 8'hE0;
            16'd21347: data <= 8'h07;
            16'd21348: data <= 8'hE0;
            16'd21349: data <= 8'h07;
            16'd21350: data <= 8'hE0;
            16'd21351: data <= 8'h07;
            16'd21352: data <= 8'hE0;
            16'd21353: data <= 8'h07;
            16'd21354: data <= 8'hE0;
            16'd21355: data <= 8'h07;
            16'd21356: data <= 8'hE0;
            16'd21357: data <= 8'h07;
            16'd21358: data <= 8'hE0;
            16'd21359: data <= 8'h07;
            16'd21360: data <= 8'hFF;
            16'd21361: data <= 8'hFF;
            16'd21362: data <= 8'hE0;
            16'd21363: data <= 8'h07;
            16'd21364: data <= 8'hE0;
            16'd21365: data <= 8'h07;
            16'd21366: data <= 8'hE0;
            16'd21367: data <= 8'h07;
            16'd21368: data <= 8'hE0;
            16'd21369: data <= 8'h07;
            16'd21370: data <= 8'hE0;
            16'd21371: data <= 8'h07;
            16'd21372: data <= 8'hE0;
            16'd21373: data <= 8'h07;
            16'd21374: data <= 8'hE0;
            16'd21375: data <= 8'h07;
            16'd21376: data <= 8'hE0;
            16'd21377: data <= 8'h07;
            16'd21378: data <= 8'hE0;
            16'd21379: data <= 8'h07;
            16'd21380: data <= 8'hE0;
            16'd21381: data <= 8'h07;
            16'd21382: data <= 8'hE0;
            16'd21383: data <= 8'h07;
            16'd21384: data <= 8'hE0;
            16'd21385: data <= 8'h07;
            16'd21386: data <= 8'hE0;
            16'd21387: data <= 8'h07;
            16'd21388: data <= 8'hE0;
            16'd21389: data <= 8'h07;
            16'd21390: data <= 8'hE0;
            16'd21391: data <= 8'h07;
            16'd21392: data <= 8'hE0;
            16'd21393: data <= 8'h07;
            16'd21394: data <= 8'hE0;
            16'd21395: data <= 8'h07;
            16'd21396: data <= 8'hE0;
            16'd21397: data <= 8'h07;
            16'd21398: data <= 8'hE0;
            16'd21399: data <= 8'h07;
            16'd21400: data <= 8'hFF;
            16'd21401: data <= 8'hFF;
            16'd21402: data <= 8'hE0;
            16'd21403: data <= 8'h07;
            16'd21404: data <= 8'hE0;
            16'd21405: data <= 8'h07;
            16'd21406: data <= 8'hE0;
            16'd21407: data <= 8'h07;
            16'd21408: data <= 8'hE0;
            16'd21409: data <= 8'h07;
            16'd21410: data <= 8'hE0;
            16'd21411: data <= 8'h07;
            16'd21412: data <= 8'hE0;
            16'd21413: data <= 8'h07;
            16'd21414: data <= 8'hE0;
            16'd21415: data <= 8'h07;
            16'd21416: data <= 8'hE0;
            16'd21417: data <= 8'h07;
            16'd21418: data <= 8'hE0;
            16'd21419: data <= 8'h07;
            16'd21420: data <= 8'hE0;
            16'd21421: data <= 8'h07;
            16'd21422: data <= 8'hE0;
            16'd21423: data <= 8'h07;
            16'd21424: data <= 8'hE0;
            16'd21425: data <= 8'h07;
            16'd21426: data <= 8'hE0;
            16'd21427: data <= 8'h07;
            16'd21428: data <= 8'hE0;
            16'd21429: data <= 8'h07;
            16'd21430: data <= 8'hE0;
            16'd21431: data <= 8'h07;
            16'd21432: data <= 8'hE0;
            16'd21433: data <= 8'h07;
            16'd21434: data <= 8'hE0;
            16'd21435: data <= 8'h07;
            16'd21436: data <= 8'hE0;
            16'd21437: data <= 8'h07;
            16'd21438: data <= 8'hE0;
            16'd21439: data <= 8'h07;
            16'd21440: data <= 8'hFF;
            16'd21441: data <= 8'hFF;
            16'd21442: data <= 8'hE0;
            16'd21443: data <= 8'h07;
            16'd21444: data <= 8'hE0;
            16'd21445: data <= 8'h07;
            16'd21446: data <= 8'hE0;
            16'd21447: data <= 8'h07;
            16'd21448: data <= 8'hE0;
            16'd21449: data <= 8'h07;
            16'd21450: data <= 8'hE0;
            16'd21451: data <= 8'h07;
            16'd21452: data <= 8'hE0;
            16'd21453: data <= 8'h07;
            16'd21454: data <= 8'hE0;
            16'd21455: data <= 8'h07;
            16'd21456: data <= 8'hE0;
            16'd21457: data <= 8'h07;
            16'd21458: data <= 8'hE0;
            16'd21459: data <= 8'h07;
            16'd21460: data <= 8'hE0;
            16'd21461: data <= 8'h07;
            16'd21462: data <= 8'hE0;
            16'd21463: data <= 8'h07;
            16'd21464: data <= 8'hE0;
            16'd21465: data <= 8'h07;
            16'd21466: data <= 8'hE0;
            16'd21467: data <= 8'h07;
            16'd21468: data <= 8'hE0;
            16'd21469: data <= 8'h07;
            16'd21470: data <= 8'hE0;
            16'd21471: data <= 8'h07;
            16'd21472: data <= 8'hE0;
            16'd21473: data <= 8'h07;
            16'd21474: data <= 8'hE0;
            16'd21475: data <= 8'h07;
            16'd21476: data <= 8'hE0;
            16'd21477: data <= 8'h07;
            16'd21478: data <= 8'hE0;
            16'd21479: data <= 8'h07;
            16'd21480: data <= 8'hFF;
            16'd21481: data <= 8'hFF;
            16'd21482: data <= 8'hE0;
            16'd21483: data <= 8'h07;
            16'd21484: data <= 8'hE0;
            16'd21485: data <= 8'h07;
            16'd21486: data <= 8'hE0;
            16'd21487: data <= 8'h07;
            16'd21488: data <= 8'hE0;
            16'd21489: data <= 8'h07;
            16'd21490: data <= 8'hE0;
            16'd21491: data <= 8'h07;
            16'd21492: data <= 8'hE0;
            16'd21493: data <= 8'h07;
            16'd21494: data <= 8'hE0;
            16'd21495: data <= 8'h07;
            16'd21496: data <= 8'hE0;
            16'd21497: data <= 8'h07;
            16'd21498: data <= 8'hE0;
            16'd21499: data <= 8'h07;
            16'd21500: data <= 8'hE0;
            16'd21501: data <= 8'h07;
            16'd21502: data <= 8'hE0;
            16'd21503: data <= 8'h07;
            16'd21504: data <= 8'hE0;
            16'd21505: data <= 8'h07;
            16'd21506: data <= 8'hE0;
            16'd21507: data <= 8'h07;
            16'd21508: data <= 8'hE0;
            16'd21509: data <= 8'h07;
            16'd21510: data <= 8'hE0;
            16'd21511: data <= 8'h07;
            16'd21512: data <= 8'hE0;
            16'd21513: data <= 8'h07;
            16'd21514: data <= 8'hE0;
            16'd21515: data <= 8'h07;
            16'd21516: data <= 8'hE0;
            16'd21517: data <= 8'h07;
            16'd21518: data <= 8'hE0;
            16'd21519: data <= 8'h07;
            16'd21520: data <= 8'hFF;
            16'd21521: data <= 8'hFF;
            16'd21522: data <= 8'hE0;
            16'd21523: data <= 8'h07;
            16'd21524: data <= 8'hE0;
            16'd21525: data <= 8'h07;
            16'd21526: data <= 8'hE0;
            16'd21527: data <= 8'h07;
            16'd21528: data <= 8'hE0;
            16'd21529: data <= 8'h07;
            16'd21530: data <= 8'hE0;
            16'd21531: data <= 8'h07;
            16'd21532: data <= 8'hE0;
            16'd21533: data <= 8'h07;
            16'd21534: data <= 8'hE0;
            16'd21535: data <= 8'h07;
            16'd21536: data <= 8'hE0;
            16'd21537: data <= 8'h07;
            16'd21538: data <= 8'hE0;
            16'd21539: data <= 8'h07;
            16'd21540: data <= 8'hE0;
            16'd21541: data <= 8'h07;
            16'd21542: data <= 8'hE0;
            16'd21543: data <= 8'h07;
            16'd21544: data <= 8'hE0;
            16'd21545: data <= 8'h07;
            16'd21546: data <= 8'hE0;
            16'd21547: data <= 8'h07;
            16'd21548: data <= 8'hE0;
            16'd21549: data <= 8'h07;
            16'd21550: data <= 8'hE0;
            16'd21551: data <= 8'h07;
            16'd21552: data <= 8'hE0;
            16'd21553: data <= 8'h07;
            16'd21554: data <= 8'hE0;
            16'd21555: data <= 8'h07;
            16'd21556: data <= 8'hE0;
            16'd21557: data <= 8'h07;
            16'd21558: data <= 8'hE0;
            16'd21559: data <= 8'h07;
            16'd21560: data <= 8'hFF;
            16'd21561: data <= 8'hFF;
            16'd21562: data <= 8'hE0;
            16'd21563: data <= 8'h07;
            16'd21564: data <= 8'hE0;
            16'd21565: data <= 8'h07;
            16'd21566: data <= 8'hE0;
            16'd21567: data <= 8'h07;
            16'd21568: data <= 8'hE0;
            16'd21569: data <= 8'h07;
            16'd21570: data <= 8'hE0;
            16'd21571: data <= 8'h07;
            16'd21572: data <= 8'hE0;
            16'd21573: data <= 8'h07;
            16'd21574: data <= 8'hE0;
            16'd21575: data <= 8'h07;
            16'd21576: data <= 8'hE0;
            16'd21577: data <= 8'h07;
            16'd21578: data <= 8'hE0;
            16'd21579: data <= 8'h07;
            16'd21580: data <= 8'hE0;
            16'd21581: data <= 8'h07;
            16'd21582: data <= 8'hE0;
            16'd21583: data <= 8'h07;
            16'd21584: data <= 8'hE0;
            16'd21585: data <= 8'h07;
            16'd21586: data <= 8'hE0;
            16'd21587: data <= 8'h07;
            16'd21588: data <= 8'hE0;
            16'd21589: data <= 8'h07;
            16'd21590: data <= 8'hE0;
            16'd21591: data <= 8'h07;
            16'd21592: data <= 8'hE0;
            16'd21593: data <= 8'h07;
            16'd21594: data <= 8'hE0;
            16'd21595: data <= 8'h07;
            16'd21596: data <= 8'hE0;
            16'd21597: data <= 8'h07;
            16'd21598: data <= 8'hE0;
            16'd21599: data <= 8'h07;
            16'd21600: data <= 8'hFF;
            16'd21601: data <= 8'hFF;
            16'd21602: data <= 8'hE0;
            16'd21603: data <= 8'h07;
            16'd21604: data <= 8'hE0;
            16'd21605: data <= 8'h07;
            16'd21606: data <= 8'hE0;
            16'd21607: data <= 8'h07;
            16'd21608: data <= 8'hE0;
            16'd21609: data <= 8'h07;
            16'd21610: data <= 8'hE0;
            16'd21611: data <= 8'h07;
            16'd21612: data <= 8'hE0;
            16'd21613: data <= 8'h07;
            16'd21614: data <= 8'hE0;
            16'd21615: data <= 8'h07;
            16'd21616: data <= 8'hE0;
            16'd21617: data <= 8'h07;
            16'd21618: data <= 8'hE0;
            16'd21619: data <= 8'h07;
            16'd21620: data <= 8'hE0;
            16'd21621: data <= 8'h07;
            16'd21622: data <= 8'hE0;
            16'd21623: data <= 8'h07;
            16'd21624: data <= 8'hE0;
            16'd21625: data <= 8'h07;
            16'd21626: data <= 8'hE0;
            16'd21627: data <= 8'h07;
            16'd21628: data <= 8'hE0;
            16'd21629: data <= 8'h07;
            16'd21630: data <= 8'hE0;
            16'd21631: data <= 8'h07;
            16'd21632: data <= 8'hE0;
            16'd21633: data <= 8'h07;
            16'd21634: data <= 8'hE0;
            16'd21635: data <= 8'h07;
            16'd21636: data <= 8'hE0;
            16'd21637: data <= 8'h07;
            16'd21638: data <= 8'hE0;
            16'd21639: data <= 8'h07;
            16'd21640: data <= 8'hFF;
            16'd21641: data <= 8'hFF;
            16'd21642: data <= 8'hE0;
            16'd21643: data <= 8'h07;
            16'd21644: data <= 8'hE0;
            16'd21645: data <= 8'h07;
            16'd21646: data <= 8'hE0;
            16'd21647: data <= 8'h07;
            16'd21648: data <= 8'hE0;
            16'd21649: data <= 8'h07;
            16'd21650: data <= 8'hE0;
            16'd21651: data <= 8'h07;
            16'd21652: data <= 8'hE0;
            16'd21653: data <= 8'h07;
            16'd21654: data <= 8'hE0;
            16'd21655: data <= 8'h07;
            16'd21656: data <= 8'hE0;
            16'd21657: data <= 8'h07;
            16'd21658: data <= 8'hE0;
            16'd21659: data <= 8'h07;
            16'd21660: data <= 8'hE0;
            16'd21661: data <= 8'h07;
            16'd21662: data <= 8'hE0;
            16'd21663: data <= 8'h07;
            16'd21664: data <= 8'hE0;
            16'd21665: data <= 8'h07;
            16'd21666: data <= 8'hE0;
            16'd21667: data <= 8'h07;
            16'd21668: data <= 8'hE0;
            16'd21669: data <= 8'h07;
            16'd21670: data <= 8'hE0;
            16'd21671: data <= 8'h07;
            16'd21672: data <= 8'hE0;
            16'd21673: data <= 8'h07;
            16'd21674: data <= 8'hE0;
            16'd21675: data <= 8'h07;
            16'd21676: data <= 8'hE0;
            16'd21677: data <= 8'h07;
            16'd21678: data <= 8'hE0;
            16'd21679: data <= 8'h07;
            16'd21680: data <= 8'hFF;
            16'd21681: data <= 8'hFF;
            16'd21682: data <= 8'hE0;
            16'd21683: data <= 8'h07;
            16'd21684: data <= 8'hE0;
            16'd21685: data <= 8'h07;
            16'd21686: data <= 8'hE0;
            16'd21687: data <= 8'h07;
            16'd21688: data <= 8'hE0;
            16'd21689: data <= 8'h07;
            16'd21690: data <= 8'hE0;
            16'd21691: data <= 8'h07;
            16'd21692: data <= 8'hE0;
            16'd21693: data <= 8'h07;
            16'd21694: data <= 8'hE0;
            16'd21695: data <= 8'h07;
            16'd21696: data <= 8'hE0;
            16'd21697: data <= 8'h07;
            16'd21698: data <= 8'hE0;
            16'd21699: data <= 8'h07;
            16'd21700: data <= 8'hE0;
            16'd21701: data <= 8'h07;
            16'd21702: data <= 8'hE0;
            16'd21703: data <= 8'h07;
            16'd21704: data <= 8'hE0;
            16'd21705: data <= 8'h07;
            16'd21706: data <= 8'hE0;
            16'd21707: data <= 8'h07;
            16'd21708: data <= 8'hE0;
            16'd21709: data <= 8'h07;
            16'd21710: data <= 8'hE0;
            16'd21711: data <= 8'h07;
            16'd21712: data <= 8'hE0;
            16'd21713: data <= 8'h07;
            16'd21714: data <= 8'hE0;
            16'd21715: data <= 8'h07;
            16'd21716: data <= 8'hE0;
            16'd21717: data <= 8'h07;
            16'd21718: data <= 8'hE0;
            16'd21719: data <= 8'h07;
            16'd21720: data <= 8'hFF;
            16'd21721: data <= 8'hFF;
            16'd21722: data <= 8'hE0;
            16'd21723: data <= 8'h07;
            16'd21724: data <= 8'hE0;
            16'd21725: data <= 8'h07;
            16'd21726: data <= 8'hE0;
            16'd21727: data <= 8'h07;
            16'd21728: data <= 8'hE0;
            16'd21729: data <= 8'h07;
            16'd21730: data <= 8'hE0;
            16'd21731: data <= 8'h07;
            16'd21732: data <= 8'hE0;
            16'd21733: data <= 8'h07;
            16'd21734: data <= 8'hE0;
            16'd21735: data <= 8'h07;
            16'd21736: data <= 8'hE0;
            16'd21737: data <= 8'h07;
            16'd21738: data <= 8'hE0;
            16'd21739: data <= 8'h07;
            16'd21740: data <= 8'hE0;
            16'd21741: data <= 8'h07;
            16'd21742: data <= 8'hE0;
            16'd21743: data <= 8'h07;
            16'd21744: data <= 8'hE0;
            16'd21745: data <= 8'h07;
            16'd21746: data <= 8'hE0;
            16'd21747: data <= 8'h07;
            16'd21748: data <= 8'hE0;
            16'd21749: data <= 8'h07;
            16'd21750: data <= 8'hE0;
            16'd21751: data <= 8'h07;
            16'd21752: data <= 8'hE0;
            16'd21753: data <= 8'h07;
            16'd21754: data <= 8'hE0;
            16'd21755: data <= 8'h07;
            16'd21756: data <= 8'hE0;
            16'd21757: data <= 8'h07;
            16'd21758: data <= 8'hE0;
            16'd21759: data <= 8'h07;
            16'd21760: data <= 8'hFF;
            16'd21761: data <= 8'hFF;
            16'd21762: data <= 8'hE0;
            16'd21763: data <= 8'h07;
            16'd21764: data <= 8'hE0;
            16'd21765: data <= 8'h07;
            16'd21766: data <= 8'hE0;
            16'd21767: data <= 8'h07;
            16'd21768: data <= 8'hE0;
            16'd21769: data <= 8'h07;
            16'd21770: data <= 8'hE0;
            16'd21771: data <= 8'h07;
            16'd21772: data <= 8'hE0;
            16'd21773: data <= 8'h07;
            16'd21774: data <= 8'hE0;
            16'd21775: data <= 8'h07;
            16'd21776: data <= 8'hE0;
            16'd21777: data <= 8'h07;
            16'd21778: data <= 8'hE0;
            16'd21779: data <= 8'h07;
            16'd21780: data <= 8'hE0;
            16'd21781: data <= 8'h07;
            16'd21782: data <= 8'hE0;
            16'd21783: data <= 8'h07;
            16'd21784: data <= 8'hE0;
            16'd21785: data <= 8'h07;
            16'd21786: data <= 8'hE0;
            16'd21787: data <= 8'h07;
            16'd21788: data <= 8'hE0;
            16'd21789: data <= 8'h07;
            16'd21790: data <= 8'hE0;
            16'd21791: data <= 8'h07;
            16'd21792: data <= 8'hE0;
            16'd21793: data <= 8'h07;
            16'd21794: data <= 8'hE0;
            16'd21795: data <= 8'h07;
            16'd21796: data <= 8'hE0;
            16'd21797: data <= 8'h07;
            16'd21798: data <= 8'hE0;
            16'd21799: data <= 8'h07;
            16'd21800: data <= 8'hFF;
            16'd21801: data <= 8'hFF;
            16'd21802: data <= 8'hE0;
            16'd21803: data <= 8'h07;
            16'd21804: data <= 8'hE0;
            16'd21805: data <= 8'h07;
            16'd21806: data <= 8'hE0;
            16'd21807: data <= 8'h07;
            16'd21808: data <= 8'hE0;
            16'd21809: data <= 8'h07;
            16'd21810: data <= 8'hE0;
            16'd21811: data <= 8'h07;
            16'd21812: data <= 8'hE0;
            16'd21813: data <= 8'h07;
            16'd21814: data <= 8'hE0;
            16'd21815: data <= 8'h07;
            16'd21816: data <= 8'hE0;
            16'd21817: data <= 8'h07;
            16'd21818: data <= 8'hE0;
            16'd21819: data <= 8'h07;
            16'd21820: data <= 8'hE0;
            16'd21821: data <= 8'h07;
            16'd21822: data <= 8'hE0;
            16'd21823: data <= 8'h07;
            16'd21824: data <= 8'hE0;
            16'd21825: data <= 8'h07;
            16'd21826: data <= 8'hE0;
            16'd21827: data <= 8'h07;
            16'd21828: data <= 8'hE0;
            16'd21829: data <= 8'h07;
            16'd21830: data <= 8'hE0;
            16'd21831: data <= 8'h07;
            16'd21832: data <= 8'hE0;
            16'd21833: data <= 8'h07;
            16'd21834: data <= 8'hE0;
            16'd21835: data <= 8'h07;
            16'd21836: data <= 8'hE0;
            16'd21837: data <= 8'h07;
            16'd21838: data <= 8'hE0;
            16'd21839: data <= 8'h07;
            16'd21840: data <= 8'hFF;
            16'd21841: data <= 8'hFF;
            16'd21842: data <= 8'hE0;
            16'd21843: data <= 8'h07;
            16'd21844: data <= 8'hE0;
            16'd21845: data <= 8'h07;
            16'd21846: data <= 8'hE0;
            16'd21847: data <= 8'h07;
            16'd21848: data <= 8'hE0;
            16'd21849: data <= 8'h07;
            16'd21850: data <= 8'hE0;
            16'd21851: data <= 8'h07;
            16'd21852: data <= 8'hE0;
            16'd21853: data <= 8'h07;
            16'd21854: data <= 8'hE0;
            16'd21855: data <= 8'h07;
            16'd21856: data <= 8'hE0;
            16'd21857: data <= 8'h07;
            16'd21858: data <= 8'hE0;
            16'd21859: data <= 8'h07;
            16'd21860: data <= 8'hE0;
            16'd21861: data <= 8'h07;
            16'd21862: data <= 8'hE0;
            16'd21863: data <= 8'h07;
            16'd21864: data <= 8'hE0;
            16'd21865: data <= 8'h07;
            16'd21866: data <= 8'hE0;
            16'd21867: data <= 8'h07;
            16'd21868: data <= 8'hE0;
            16'd21869: data <= 8'h07;
            16'd21870: data <= 8'hE0;
            16'd21871: data <= 8'h07;
            16'd21872: data <= 8'hE0;
            16'd21873: data <= 8'h07;
            16'd21874: data <= 8'hE0;
            16'd21875: data <= 8'h07;
            16'd21876: data <= 8'hE0;
            16'd21877: data <= 8'h07;
            16'd21878: data <= 8'hE0;
            16'd21879: data <= 8'h07;
            16'd21880: data <= 8'hFF;
            16'd21881: data <= 8'hFF;
            16'd21882: data <= 8'hE0;
            16'd21883: data <= 8'h07;
            16'd21884: data <= 8'hE0;
            16'd21885: data <= 8'h07;
            16'd21886: data <= 8'hE0;
            16'd21887: data <= 8'h07;
            16'd21888: data <= 8'hE0;
            16'd21889: data <= 8'h07;
            16'd21890: data <= 8'hE0;
            16'd21891: data <= 8'h07;
            16'd21892: data <= 8'hE0;
            16'd21893: data <= 8'h07;
            16'd21894: data <= 8'hE0;
            16'd21895: data <= 8'h07;
            16'd21896: data <= 8'hE0;
            16'd21897: data <= 8'h07;
            16'd21898: data <= 8'hE0;
            16'd21899: data <= 8'h07;
            16'd21900: data <= 8'hE0;
            16'd21901: data <= 8'h07;
            16'd21902: data <= 8'hE0;
            16'd21903: data <= 8'h07;
            16'd21904: data <= 8'hE0;
            16'd21905: data <= 8'h07;
            16'd21906: data <= 8'hE0;
            16'd21907: data <= 8'h07;
            16'd21908: data <= 8'hE0;
            16'd21909: data <= 8'h07;
            16'd21910: data <= 8'hE0;
            16'd21911: data <= 8'h07;
            16'd21912: data <= 8'hE0;
            16'd21913: data <= 8'h07;
            16'd21914: data <= 8'hE0;
            16'd21915: data <= 8'h07;
            16'd21916: data <= 8'hE0;
            16'd21917: data <= 8'h07;
            16'd21918: data <= 8'hE0;
            16'd21919: data <= 8'h07;
            16'd21920: data <= 8'hFF;
            16'd21921: data <= 8'hFF;
            16'd21922: data <= 8'hE0;
            16'd21923: data <= 8'h07;
            16'd21924: data <= 8'hE0;
            16'd21925: data <= 8'h07;
            16'd21926: data <= 8'hE0;
            16'd21927: data <= 8'h07;
            16'd21928: data <= 8'hE0;
            16'd21929: data <= 8'h07;
            16'd21930: data <= 8'hE0;
            16'd21931: data <= 8'h07;
            16'd21932: data <= 8'hE0;
            16'd21933: data <= 8'h07;
            16'd21934: data <= 8'hE0;
            16'd21935: data <= 8'h07;
            16'd21936: data <= 8'hE0;
            16'd21937: data <= 8'h07;
            16'd21938: data <= 8'hE0;
            16'd21939: data <= 8'h07;
            16'd21940: data <= 8'hE0;
            16'd21941: data <= 8'h07;
            16'd21942: data <= 8'hE0;
            16'd21943: data <= 8'h07;
            16'd21944: data <= 8'hE0;
            16'd21945: data <= 8'h07;
            16'd21946: data <= 8'hE0;
            16'd21947: data <= 8'h07;
            16'd21948: data <= 8'hE0;
            16'd21949: data <= 8'h07;
            16'd21950: data <= 8'hE0;
            16'd21951: data <= 8'h07;
            16'd21952: data <= 8'hE0;
            16'd21953: data <= 8'h07;
            16'd21954: data <= 8'hE0;
            16'd21955: data <= 8'h07;
            16'd21956: data <= 8'hE0;
            16'd21957: data <= 8'h07;
            16'd21958: data <= 8'hE0;
            16'd21959: data <= 8'h07;
            16'd21960: data <= 8'hFF;
            16'd21961: data <= 8'hFF;
            16'd21962: data <= 8'hE0;
            16'd21963: data <= 8'h07;
            16'd21964: data <= 8'hE0;
            16'd21965: data <= 8'h07;
            16'd21966: data <= 8'hE0;
            16'd21967: data <= 8'h07;
            16'd21968: data <= 8'hE0;
            16'd21969: data <= 8'h07;
            16'd21970: data <= 8'hE0;
            16'd21971: data <= 8'h07;
            16'd21972: data <= 8'hE0;
            16'd21973: data <= 8'h07;
            16'd21974: data <= 8'hE0;
            16'd21975: data <= 8'h07;
            16'd21976: data <= 8'hE0;
            16'd21977: data <= 8'h07;
            16'd21978: data <= 8'hE0;
            16'd21979: data <= 8'h07;
            16'd21980: data <= 8'hE0;
            16'd21981: data <= 8'h07;
            16'd21982: data <= 8'hE0;
            16'd21983: data <= 8'h07;
            16'd21984: data <= 8'hE0;
            16'd21985: data <= 8'h07;
            16'd21986: data <= 8'hE0;
            16'd21987: data <= 8'h07;
            16'd21988: data <= 8'hE0;
            16'd21989: data <= 8'h07;
            16'd21990: data <= 8'hE0;
            16'd21991: data <= 8'h07;
            16'd21992: data <= 8'hE0;
            16'd21993: data <= 8'h07;
            16'd21994: data <= 8'hE0;
            16'd21995: data <= 8'h07;
            16'd21996: data <= 8'hE0;
            16'd21997: data <= 8'h07;
            16'd21998: data <= 8'hE0;
            16'd21999: data <= 8'h07;
            16'd22000: data <= 8'hFF;
            16'd22001: data <= 8'hFF;
            16'd22002: data <= 8'hE0;
            16'd22003: data <= 8'h07;
            16'd22004: data <= 8'hE0;
            16'd22005: data <= 8'h07;
            16'd22006: data <= 8'hE0;
            16'd22007: data <= 8'h07;
            16'd22008: data <= 8'hE0;
            16'd22009: data <= 8'h07;
            16'd22010: data <= 8'hE0;
            16'd22011: data <= 8'h07;
            16'd22012: data <= 8'hE0;
            16'd22013: data <= 8'h07;
            16'd22014: data <= 8'hE0;
            16'd22015: data <= 8'h07;
            16'd22016: data <= 8'hE0;
            16'd22017: data <= 8'h07;
            16'd22018: data <= 8'hE0;
            16'd22019: data <= 8'h07;
            16'd22020: data <= 8'hE0;
            16'd22021: data <= 8'h07;
            16'd22022: data <= 8'hE0;
            16'd22023: data <= 8'h07;
            16'd22024: data <= 8'hE0;
            16'd22025: data <= 8'h07;
            16'd22026: data <= 8'hE0;
            16'd22027: data <= 8'h07;
            16'd22028: data <= 8'hE0;
            16'd22029: data <= 8'h07;
            16'd22030: data <= 8'hE0;
            16'd22031: data <= 8'h07;
            16'd22032: data <= 8'hE0;
            16'd22033: data <= 8'h07;
            16'd22034: data <= 8'hE0;
            16'd22035: data <= 8'h07;
            16'd22036: data <= 8'hE0;
            16'd22037: data <= 8'h07;
            16'd22038: data <= 8'hE0;
            16'd22039: data <= 8'h07;
            16'd22040: data <= 8'hFF;
            16'd22041: data <= 8'hFF;
            16'd22042: data <= 8'hE0;
            16'd22043: data <= 8'h07;
            16'd22044: data <= 8'hE0;
            16'd22045: data <= 8'h07;
            16'd22046: data <= 8'hE0;
            16'd22047: data <= 8'h07;
            16'd22048: data <= 8'hE0;
            16'd22049: data <= 8'h07;
            16'd22050: data <= 8'hE0;
            16'd22051: data <= 8'h07;
            16'd22052: data <= 8'hE0;
            16'd22053: data <= 8'h07;
            16'd22054: data <= 8'hE0;
            16'd22055: data <= 8'h07;
            16'd22056: data <= 8'hE0;
            16'd22057: data <= 8'h07;
            16'd22058: data <= 8'hE0;
            16'd22059: data <= 8'h07;
            16'd22060: data <= 8'hE0;
            16'd22061: data <= 8'h07;
            16'd22062: data <= 8'hE0;
            16'd22063: data <= 8'h07;
            16'd22064: data <= 8'hE0;
            16'd22065: data <= 8'h07;
            16'd22066: data <= 8'hE0;
            16'd22067: data <= 8'h07;
            16'd22068: data <= 8'hE0;
            16'd22069: data <= 8'h07;
            16'd22070: data <= 8'hE0;
            16'd22071: data <= 8'h07;
            16'd22072: data <= 8'hE0;
            16'd22073: data <= 8'h07;
            16'd22074: data <= 8'hE0;
            16'd22075: data <= 8'h07;
            16'd22076: data <= 8'hE0;
            16'd22077: data <= 8'h07;
            16'd22078: data <= 8'hE0;
            16'd22079: data <= 8'h07;
            16'd22080: data <= 8'hFF;
            16'd22081: data <= 8'hFF;
            16'd22082: data <= 8'hE0;
            16'd22083: data <= 8'h07;
            16'd22084: data <= 8'hE0;
            16'd22085: data <= 8'h07;
            16'd22086: data <= 8'hE0;
            16'd22087: data <= 8'h07;
            16'd22088: data <= 8'hE0;
            16'd22089: data <= 8'h07;
            16'd22090: data <= 8'hE0;
            16'd22091: data <= 8'h07;
            16'd22092: data <= 8'hE0;
            16'd22093: data <= 8'h07;
            16'd22094: data <= 8'hE0;
            16'd22095: data <= 8'h07;
            16'd22096: data <= 8'hE0;
            16'd22097: data <= 8'h07;
            16'd22098: data <= 8'hE0;
            16'd22099: data <= 8'h07;
            16'd22100: data <= 8'hE0;
            16'd22101: data <= 8'h07;
            16'd22102: data <= 8'hE0;
            16'd22103: data <= 8'h07;
            16'd22104: data <= 8'hE0;
            16'd22105: data <= 8'h07;
            16'd22106: data <= 8'hE0;
            16'd22107: data <= 8'h07;
            16'd22108: data <= 8'hE0;
            16'd22109: data <= 8'h07;
            16'd22110: data <= 8'hE0;
            16'd22111: data <= 8'h07;
            16'd22112: data <= 8'hE0;
            16'd22113: data <= 8'h07;
            16'd22114: data <= 8'hE0;
            16'd22115: data <= 8'h07;
            16'd22116: data <= 8'hE0;
            16'd22117: data <= 8'h07;
            16'd22118: data <= 8'hE0;
            16'd22119: data <= 8'h07;
            16'd22120: data <= 8'hFF;
            16'd22121: data <= 8'hFF;
            16'd22122: data <= 8'hE0;
            16'd22123: data <= 8'h07;
            16'd22124: data <= 8'hE0;
            16'd22125: data <= 8'h07;
            16'd22126: data <= 8'hE0;
            16'd22127: data <= 8'h07;
            16'd22128: data <= 8'hE0;
            16'd22129: data <= 8'h07;
            16'd22130: data <= 8'hE0;
            16'd22131: data <= 8'h07;
            16'd22132: data <= 8'hE0;
            16'd22133: data <= 8'h07;
            16'd22134: data <= 8'hE0;
            16'd22135: data <= 8'h07;
            16'd22136: data <= 8'hE0;
            16'd22137: data <= 8'h07;
            16'd22138: data <= 8'hE0;
            16'd22139: data <= 8'h07;
            16'd22140: data <= 8'hE0;
            16'd22141: data <= 8'h07;
            16'd22142: data <= 8'hE0;
            16'd22143: data <= 8'h07;
            16'd22144: data <= 8'hE0;
            16'd22145: data <= 8'h07;
            16'd22146: data <= 8'hE0;
            16'd22147: data <= 8'h07;
            16'd22148: data <= 8'hE0;
            16'd22149: data <= 8'h07;
            16'd22150: data <= 8'hE0;
            16'd22151: data <= 8'h07;
            16'd22152: data <= 8'hE0;
            16'd22153: data <= 8'h07;
            16'd22154: data <= 8'hE0;
            16'd22155: data <= 8'h07;
            16'd22156: data <= 8'hE0;
            16'd22157: data <= 8'h07;
            16'd22158: data <= 8'hE0;
            16'd22159: data <= 8'h07;
            16'd22160: data <= 8'hFF;
            16'd22161: data <= 8'hFF;
            16'd22162: data <= 8'hE0;
            16'd22163: data <= 8'h07;
            16'd22164: data <= 8'hE0;
            16'd22165: data <= 8'h07;
            16'd22166: data <= 8'hE0;
            16'd22167: data <= 8'h07;
            16'd22168: data <= 8'hE0;
            16'd22169: data <= 8'h07;
            16'd22170: data <= 8'hE0;
            16'd22171: data <= 8'h07;
            16'd22172: data <= 8'hE0;
            16'd22173: data <= 8'h07;
            16'd22174: data <= 8'hE0;
            16'd22175: data <= 8'h07;
            16'd22176: data <= 8'hE0;
            16'd22177: data <= 8'h07;
            16'd22178: data <= 8'hE0;
            16'd22179: data <= 8'h07;
            16'd22180: data <= 8'hE0;
            16'd22181: data <= 8'h07;
            16'd22182: data <= 8'hE0;
            16'd22183: data <= 8'h07;
            16'd22184: data <= 8'hE0;
            16'd22185: data <= 8'h07;
            16'd22186: data <= 8'hE0;
            16'd22187: data <= 8'h07;
            16'd22188: data <= 8'hE0;
            16'd22189: data <= 8'h07;
            16'd22190: data <= 8'hE0;
            16'd22191: data <= 8'h07;
            16'd22192: data <= 8'hE0;
            16'd22193: data <= 8'h07;
            16'd22194: data <= 8'hE0;
            16'd22195: data <= 8'h07;
            16'd22196: data <= 8'hE0;
            16'd22197: data <= 8'h07;
            16'd22198: data <= 8'hE0;
            16'd22199: data <= 8'h07;
            16'd22200: data <= 8'hFF;
            16'd22201: data <= 8'hFF;
            16'd22202: data <= 8'hE0;
            16'd22203: data <= 8'h07;
            16'd22204: data <= 8'hE0;
            16'd22205: data <= 8'h07;
            16'd22206: data <= 8'hE0;
            16'd22207: data <= 8'h07;
            16'd22208: data <= 8'hE0;
            16'd22209: data <= 8'h07;
            16'd22210: data <= 8'hE0;
            16'd22211: data <= 8'h07;
            16'd22212: data <= 8'hE0;
            16'd22213: data <= 8'h07;
            16'd22214: data <= 8'hE0;
            16'd22215: data <= 8'h07;
            16'd22216: data <= 8'hE0;
            16'd22217: data <= 8'h07;
            16'd22218: data <= 8'hE0;
            16'd22219: data <= 8'h07;
            16'd22220: data <= 8'hE0;
            16'd22221: data <= 8'h07;
            16'd22222: data <= 8'hE0;
            16'd22223: data <= 8'h07;
            16'd22224: data <= 8'hE0;
            16'd22225: data <= 8'h07;
            16'd22226: data <= 8'hE0;
            16'd22227: data <= 8'h07;
            16'd22228: data <= 8'hE0;
            16'd22229: data <= 8'h07;
            16'd22230: data <= 8'hE0;
            16'd22231: data <= 8'h07;
            16'd22232: data <= 8'hE0;
            16'd22233: data <= 8'h07;
            16'd22234: data <= 8'hE0;
            16'd22235: data <= 8'h07;
            16'd22236: data <= 8'hE0;
            16'd22237: data <= 8'h07;
            16'd22238: data <= 8'hE0;
            16'd22239: data <= 8'h07;
            16'd22240: data <= 8'hFF;
            16'd22241: data <= 8'hFF;
            16'd22242: data <= 8'hE0;
            16'd22243: data <= 8'h07;
            16'd22244: data <= 8'hE0;
            16'd22245: data <= 8'h07;
            16'd22246: data <= 8'hE0;
            16'd22247: data <= 8'h07;
            16'd22248: data <= 8'hE0;
            16'd22249: data <= 8'h07;
            16'd22250: data <= 8'hE0;
            16'd22251: data <= 8'h07;
            16'd22252: data <= 8'hE0;
            16'd22253: data <= 8'h07;
            16'd22254: data <= 8'hE0;
            16'd22255: data <= 8'h07;
            16'd22256: data <= 8'hE0;
            16'd22257: data <= 8'h07;
            16'd22258: data <= 8'hE0;
            16'd22259: data <= 8'h07;
            16'd22260: data <= 8'hE0;
            16'd22261: data <= 8'h07;
            16'd22262: data <= 8'hE0;
            16'd22263: data <= 8'h07;
            16'd22264: data <= 8'hE0;
            16'd22265: data <= 8'h07;
            16'd22266: data <= 8'hE0;
            16'd22267: data <= 8'h07;
            16'd22268: data <= 8'hE0;
            16'd22269: data <= 8'h07;
            16'd22270: data <= 8'hE0;
            16'd22271: data <= 8'h07;
            16'd22272: data <= 8'hE0;
            16'd22273: data <= 8'h07;
            16'd22274: data <= 8'hE0;
            16'd22275: data <= 8'h07;
            16'd22276: data <= 8'hE0;
            16'd22277: data <= 8'h07;
            16'd22278: data <= 8'hE0;
            16'd22279: data <= 8'h07;
            16'd22280: data <= 8'hFF;
            16'd22281: data <= 8'hFF;
            16'd22282: data <= 8'hE0;
            16'd22283: data <= 8'h07;
            16'd22284: data <= 8'hE0;
            16'd22285: data <= 8'h07;
            16'd22286: data <= 8'hE0;
            16'd22287: data <= 8'h07;
            16'd22288: data <= 8'hE0;
            16'd22289: data <= 8'h07;
            16'd22290: data <= 8'hE0;
            16'd22291: data <= 8'h07;
            16'd22292: data <= 8'hE0;
            16'd22293: data <= 8'h07;
            16'd22294: data <= 8'hE0;
            16'd22295: data <= 8'h07;
            16'd22296: data <= 8'hE0;
            16'd22297: data <= 8'h07;
            16'd22298: data <= 8'hE0;
            16'd22299: data <= 8'h07;
            16'd22300: data <= 8'hE0;
            16'd22301: data <= 8'h07;
            16'd22302: data <= 8'hE0;
            16'd22303: data <= 8'h07;
            16'd22304: data <= 8'hE0;
            16'd22305: data <= 8'h07;
            16'd22306: data <= 8'hE0;
            16'd22307: data <= 8'h07;
            16'd22308: data <= 8'hE0;
            16'd22309: data <= 8'h07;
            16'd22310: data <= 8'hE0;
            16'd22311: data <= 8'h07;
            16'd22312: data <= 8'hE0;
            16'd22313: data <= 8'h07;
            16'd22314: data <= 8'hE0;
            16'd22315: data <= 8'h07;
            16'd22316: data <= 8'hE0;
            16'd22317: data <= 8'h07;
            16'd22318: data <= 8'hE0;
            16'd22319: data <= 8'h07;
            16'd22320: data <= 8'hFF;
            16'd22321: data <= 8'hFF;
            16'd22322: data <= 8'hE0;
            16'd22323: data <= 8'h07;
            16'd22324: data <= 8'hE0;
            16'd22325: data <= 8'h07;
            16'd22326: data <= 8'hE0;
            16'd22327: data <= 8'h07;
            16'd22328: data <= 8'hE0;
            16'd22329: data <= 8'h07;
            16'd22330: data <= 8'hE0;
            16'd22331: data <= 8'h07;
            16'd22332: data <= 8'hE0;
            16'd22333: data <= 8'h07;
            16'd22334: data <= 8'hE0;
            16'd22335: data <= 8'h07;
            16'd22336: data <= 8'hE0;
            16'd22337: data <= 8'h07;
            16'd22338: data <= 8'hE0;
            16'd22339: data <= 8'h07;
            16'd22340: data <= 8'hE0;
            16'd22341: data <= 8'h07;
            16'd22342: data <= 8'hE0;
            16'd22343: data <= 8'h07;
            16'd22344: data <= 8'hE0;
            16'd22345: data <= 8'h07;
            16'd22346: data <= 8'hE0;
            16'd22347: data <= 8'h07;
            16'd22348: data <= 8'hE0;
            16'd22349: data <= 8'h07;
            16'd22350: data <= 8'hE0;
            16'd22351: data <= 8'h07;
            16'd22352: data <= 8'hE0;
            16'd22353: data <= 8'h07;
            16'd22354: data <= 8'hE0;
            16'd22355: data <= 8'h07;
            16'd22356: data <= 8'hE0;
            16'd22357: data <= 8'h07;
            16'd22358: data <= 8'hE0;
            16'd22359: data <= 8'h07;
            16'd22360: data <= 8'hFF;
            16'd22361: data <= 8'hFF;
            16'd22362: data <= 8'hE0;
            16'd22363: data <= 8'h07;
            16'd22364: data <= 8'hE0;
            16'd22365: data <= 8'h07;
            16'd22366: data <= 8'hE0;
            16'd22367: data <= 8'h07;
            16'd22368: data <= 8'hE0;
            16'd22369: data <= 8'h07;
            16'd22370: data <= 8'hE0;
            16'd22371: data <= 8'h07;
            16'd22372: data <= 8'hE0;
            16'd22373: data <= 8'h07;
            16'd22374: data <= 8'hE0;
            16'd22375: data <= 8'h07;
            16'd22376: data <= 8'hE0;
            16'd22377: data <= 8'h07;
            16'd22378: data <= 8'hE0;
            16'd22379: data <= 8'h07;
            16'd22380: data <= 8'hE0;
            16'd22381: data <= 8'h07;
            16'd22382: data <= 8'hE0;
            16'd22383: data <= 8'h07;
            16'd22384: data <= 8'hE0;
            16'd22385: data <= 8'h07;
            16'd22386: data <= 8'hE0;
            16'd22387: data <= 8'h07;
            16'd22388: data <= 8'hE0;
            16'd22389: data <= 8'h07;
            16'd22390: data <= 8'hE0;
            16'd22391: data <= 8'h07;
            16'd22392: data <= 8'hE0;
            16'd22393: data <= 8'h07;
            16'd22394: data <= 8'hE0;
            16'd22395: data <= 8'h07;
            16'd22396: data <= 8'hE0;
            16'd22397: data <= 8'h07;
            16'd22398: data <= 8'hE0;
            16'd22399: data <= 8'h07;
            16'd22400: data <= 8'hFF;
            16'd22401: data <= 8'hFF;
            16'd22402: data <= 8'hE0;
            16'd22403: data <= 8'h07;
            16'd22404: data <= 8'hE0;
            16'd22405: data <= 8'h07;
            16'd22406: data <= 8'hE0;
            16'd22407: data <= 8'h07;
            16'd22408: data <= 8'hE0;
            16'd22409: data <= 8'h07;
            16'd22410: data <= 8'hE0;
            16'd22411: data <= 8'h07;
            16'd22412: data <= 8'hE0;
            16'd22413: data <= 8'h07;
            16'd22414: data <= 8'hE0;
            16'd22415: data <= 8'h07;
            16'd22416: data <= 8'hE0;
            16'd22417: data <= 8'h07;
            16'd22418: data <= 8'hE0;
            16'd22419: data <= 8'h07;
            16'd22420: data <= 8'hE0;
            16'd22421: data <= 8'h07;
            16'd22422: data <= 8'hE0;
            16'd22423: data <= 8'h07;
            16'd22424: data <= 8'hE0;
            16'd22425: data <= 8'h07;
            16'd22426: data <= 8'hE0;
            16'd22427: data <= 8'h07;
            16'd22428: data <= 8'hE0;
            16'd22429: data <= 8'h07;
            16'd22430: data <= 8'hE0;
            16'd22431: data <= 8'h07;
            16'd22432: data <= 8'hE0;
            16'd22433: data <= 8'h07;
            16'd22434: data <= 8'hE0;
            16'd22435: data <= 8'h07;
            16'd22436: data <= 8'hE0;
            16'd22437: data <= 8'h07;
            16'd22438: data <= 8'hE0;
            16'd22439: data <= 8'h07;
            16'd22440: data <= 8'hFF;
            16'd22441: data <= 8'hFF;
            16'd22442: data <= 8'hE0;
            16'd22443: data <= 8'h07;
            16'd22444: data <= 8'hE0;
            16'd22445: data <= 8'h07;
            16'd22446: data <= 8'hE0;
            16'd22447: data <= 8'h07;
            16'd22448: data <= 8'hE0;
            16'd22449: data <= 8'h07;
            16'd22450: data <= 8'hE0;
            16'd22451: data <= 8'h07;
            16'd22452: data <= 8'hE0;
            16'd22453: data <= 8'h07;
            16'd22454: data <= 8'hE0;
            16'd22455: data <= 8'h07;
            16'd22456: data <= 8'hE0;
            16'd22457: data <= 8'h07;
            16'd22458: data <= 8'hE0;
            16'd22459: data <= 8'h07;
            16'd22460: data <= 8'hE0;
            16'd22461: data <= 8'h07;
            16'd22462: data <= 8'hE0;
            16'd22463: data <= 8'h07;
            16'd22464: data <= 8'hE0;
            16'd22465: data <= 8'h07;
            16'd22466: data <= 8'hE0;
            16'd22467: data <= 8'h07;
            16'd22468: data <= 8'hE0;
            16'd22469: data <= 8'h07;
            16'd22470: data <= 8'hE0;
            16'd22471: data <= 8'h07;
            16'd22472: data <= 8'hE0;
            16'd22473: data <= 8'h07;
            16'd22474: data <= 8'hE0;
            16'd22475: data <= 8'h07;
            16'd22476: data <= 8'hE0;
            16'd22477: data <= 8'h07;
            16'd22478: data <= 8'hE0;
            16'd22479: data <= 8'h07;
            16'd22480: data <= 8'hFF;
            16'd22481: data <= 8'hFF;
            16'd22482: data <= 8'hE0;
            16'd22483: data <= 8'h07;
            16'd22484: data <= 8'hE0;
            16'd22485: data <= 8'h07;
            16'd22486: data <= 8'hE0;
            16'd22487: data <= 8'h07;
            16'd22488: data <= 8'hE0;
            16'd22489: data <= 8'h07;
            16'd22490: data <= 8'hE0;
            16'd22491: data <= 8'h07;
            16'd22492: data <= 8'hE0;
            16'd22493: data <= 8'h07;
            16'd22494: data <= 8'hE0;
            16'd22495: data <= 8'h07;
            16'd22496: data <= 8'hE0;
            16'd22497: data <= 8'h07;
            16'd22498: data <= 8'hE0;
            16'd22499: data <= 8'h07;
            16'd22500: data <= 8'hE0;
            16'd22501: data <= 8'h07;
            16'd22502: data <= 8'hE0;
            16'd22503: data <= 8'h07;
            16'd22504: data <= 8'hE0;
            16'd22505: data <= 8'h07;
            16'd22506: data <= 8'hE0;
            16'd22507: data <= 8'h07;
            16'd22508: data <= 8'hE0;
            16'd22509: data <= 8'h07;
            16'd22510: data <= 8'hE0;
            16'd22511: data <= 8'h07;
            16'd22512: data <= 8'hE0;
            16'd22513: data <= 8'h07;
            16'd22514: data <= 8'hE0;
            16'd22515: data <= 8'h07;
            16'd22516: data <= 8'hE0;
            16'd22517: data <= 8'h07;
            16'd22518: data <= 8'hE0;
            16'd22519: data <= 8'h07;
            16'd22520: data <= 8'hFF;
            16'd22521: data <= 8'hFF;
            16'd22522: data <= 8'hE0;
            16'd22523: data <= 8'h07;
            16'd22524: data <= 8'hE0;
            16'd22525: data <= 8'h07;
            16'd22526: data <= 8'hE0;
            16'd22527: data <= 8'h07;
            16'd22528: data <= 8'hE0;
            16'd22529: data <= 8'h07;
            16'd22530: data <= 8'hE0;
            16'd22531: data <= 8'h07;
            16'd22532: data <= 8'hE0;
            16'd22533: data <= 8'h07;
            16'd22534: data <= 8'hE0;
            16'd22535: data <= 8'h07;
            16'd22536: data <= 8'hE0;
            16'd22537: data <= 8'h07;
            16'd22538: data <= 8'hE0;
            16'd22539: data <= 8'h07;
            16'd22540: data <= 8'hE0;
            16'd22541: data <= 8'h07;
            16'd22542: data <= 8'hE0;
            16'd22543: data <= 8'h07;
            16'd22544: data <= 8'hE0;
            16'd22545: data <= 8'h07;
            16'd22546: data <= 8'hE0;
            16'd22547: data <= 8'h07;
            16'd22548: data <= 8'hE0;
            16'd22549: data <= 8'h07;
            16'd22550: data <= 8'hE0;
            16'd22551: data <= 8'h07;
            16'd22552: data <= 8'hE0;
            16'd22553: data <= 8'h07;
            16'd22554: data <= 8'hE0;
            16'd22555: data <= 8'h07;
            16'd22556: data <= 8'hE0;
            16'd22557: data <= 8'h07;
            16'd22558: data <= 8'hE0;
            16'd22559: data <= 8'h07;
            16'd22560: data <= 8'hFF;
            16'd22561: data <= 8'hFF;
            16'd22562: data <= 8'hE0;
            16'd22563: data <= 8'h07;
            16'd22564: data <= 8'hE0;
            16'd22565: data <= 8'h07;
            16'd22566: data <= 8'hE0;
            16'd22567: data <= 8'h07;
            16'd22568: data <= 8'hE0;
            16'd22569: data <= 8'h07;
            16'd22570: data <= 8'hE0;
            16'd22571: data <= 8'h07;
            16'd22572: data <= 8'hE0;
            16'd22573: data <= 8'h07;
            16'd22574: data <= 8'hE0;
            16'd22575: data <= 8'h07;
            16'd22576: data <= 8'hE0;
            16'd22577: data <= 8'h07;
            16'd22578: data <= 8'hE0;
            16'd22579: data <= 8'h07;
            16'd22580: data <= 8'hE0;
            16'd22581: data <= 8'h07;
            16'd22582: data <= 8'hE0;
            16'd22583: data <= 8'h07;
            16'd22584: data <= 8'hE0;
            16'd22585: data <= 8'h07;
            16'd22586: data <= 8'hE0;
            16'd22587: data <= 8'h07;
            16'd22588: data <= 8'hE0;
            16'd22589: data <= 8'h07;
            16'd22590: data <= 8'hE0;
            16'd22591: data <= 8'h07;
            16'd22592: data <= 8'hE0;
            16'd22593: data <= 8'h07;
            16'd22594: data <= 8'hE0;
            16'd22595: data <= 8'h07;
            16'd22596: data <= 8'hE0;
            16'd22597: data <= 8'h07;
            16'd22598: data <= 8'hE0;
            16'd22599: data <= 8'h07;
            16'd22600: data <= 8'hFF;
            16'd22601: data <= 8'hFF;
            16'd22602: data <= 8'hE0;
            16'd22603: data <= 8'h07;
            16'd22604: data <= 8'hE0;
            16'd22605: data <= 8'h07;
            16'd22606: data <= 8'hE0;
            16'd22607: data <= 8'h07;
            16'd22608: data <= 8'hE0;
            16'd22609: data <= 8'h07;
            16'd22610: data <= 8'hE0;
            16'd22611: data <= 8'h07;
            16'd22612: data <= 8'hE0;
            16'd22613: data <= 8'h07;
            16'd22614: data <= 8'hE0;
            16'd22615: data <= 8'h07;
            16'd22616: data <= 8'hE0;
            16'd22617: data <= 8'h07;
            16'd22618: data <= 8'hE0;
            16'd22619: data <= 8'h07;
            16'd22620: data <= 8'hE0;
            16'd22621: data <= 8'h07;
            16'd22622: data <= 8'hE0;
            16'd22623: data <= 8'h07;
            16'd22624: data <= 8'hE0;
            16'd22625: data <= 8'h07;
            16'd22626: data <= 8'hE0;
            16'd22627: data <= 8'h07;
            16'd22628: data <= 8'hE0;
            16'd22629: data <= 8'h07;
            16'd22630: data <= 8'hE0;
            16'd22631: data <= 8'h07;
            16'd22632: data <= 8'hE0;
            16'd22633: data <= 8'h07;
            16'd22634: data <= 8'hE0;
            16'd22635: data <= 8'h07;
            16'd22636: data <= 8'hE0;
            16'd22637: data <= 8'h07;
            16'd22638: data <= 8'hE0;
            16'd22639: data <= 8'h07;
            16'd22640: data <= 8'hFF;
            16'd22641: data <= 8'hFF;
            16'd22642: data <= 8'hE0;
            16'd22643: data <= 8'h07;
            16'd22644: data <= 8'hE0;
            16'd22645: data <= 8'h07;
            16'd22646: data <= 8'hE0;
            16'd22647: data <= 8'h07;
            16'd22648: data <= 8'hE0;
            16'd22649: data <= 8'h07;
            16'd22650: data <= 8'hE0;
            16'd22651: data <= 8'h07;
            16'd22652: data <= 8'hE0;
            16'd22653: data <= 8'h07;
            16'd22654: data <= 8'hE0;
            16'd22655: data <= 8'h07;
            16'd22656: data <= 8'hE0;
            16'd22657: data <= 8'h07;
            16'd22658: data <= 8'hE0;
            16'd22659: data <= 8'h07;
            16'd22660: data <= 8'hE0;
            16'd22661: data <= 8'h07;
            16'd22662: data <= 8'hE0;
            16'd22663: data <= 8'h07;
            16'd22664: data <= 8'hE0;
            16'd22665: data <= 8'h07;
            16'd22666: data <= 8'hE0;
            16'd22667: data <= 8'h07;
            16'd22668: data <= 8'hE0;
            16'd22669: data <= 8'h07;
            16'd22670: data <= 8'hE0;
            16'd22671: data <= 8'h07;
            16'd22672: data <= 8'hE0;
            16'd22673: data <= 8'h07;
            16'd22674: data <= 8'hE0;
            16'd22675: data <= 8'h07;
            16'd22676: data <= 8'hE0;
            16'd22677: data <= 8'h07;
            16'd22678: data <= 8'hE0;
            16'd22679: data <= 8'h07;
            16'd22680: data <= 8'hFF;
            16'd22681: data <= 8'hFF;
            16'd22682: data <= 8'hE0;
            16'd22683: data <= 8'h07;
            16'd22684: data <= 8'hE0;
            16'd22685: data <= 8'h07;
            16'd22686: data <= 8'hE0;
            16'd22687: data <= 8'h07;
            16'd22688: data <= 8'hE0;
            16'd22689: data <= 8'h07;
            16'd22690: data <= 8'hE0;
            16'd22691: data <= 8'h07;
            16'd22692: data <= 8'hE0;
            16'd22693: data <= 8'h07;
            16'd22694: data <= 8'hE0;
            16'd22695: data <= 8'h07;
            16'd22696: data <= 8'hE0;
            16'd22697: data <= 8'h07;
            16'd22698: data <= 8'hE0;
            16'd22699: data <= 8'h07;
            16'd22700: data <= 8'hE0;
            16'd22701: data <= 8'h07;
            16'd22702: data <= 8'hE0;
            16'd22703: data <= 8'h07;
            16'd22704: data <= 8'hE0;
            16'd22705: data <= 8'h07;
            16'd22706: data <= 8'hE0;
            16'd22707: data <= 8'h07;
            16'd22708: data <= 8'hE0;
            16'd22709: data <= 8'h07;
            16'd22710: data <= 8'hE0;
            16'd22711: data <= 8'h07;
            16'd22712: data <= 8'hE0;
            16'd22713: data <= 8'h07;
            16'd22714: data <= 8'hE0;
            16'd22715: data <= 8'h07;
            16'd22716: data <= 8'hE0;
            16'd22717: data <= 8'h07;
            16'd22718: data <= 8'hE0;
            16'd22719: data <= 8'h07;
            16'd22720: data <= 8'hFF;
            16'd22721: data <= 8'hFF;
            16'd22722: data <= 8'hE0;
            16'd22723: data <= 8'h07;
            16'd22724: data <= 8'hE0;
            16'd22725: data <= 8'h07;
            16'd22726: data <= 8'hE0;
            16'd22727: data <= 8'h07;
            16'd22728: data <= 8'hE0;
            16'd22729: data <= 8'h07;
            16'd22730: data <= 8'hE0;
            16'd22731: data <= 8'h07;
            16'd22732: data <= 8'hE0;
            16'd22733: data <= 8'h07;
            16'd22734: data <= 8'hE0;
            16'd22735: data <= 8'h07;
            16'd22736: data <= 8'hE0;
            16'd22737: data <= 8'h07;
            16'd22738: data <= 8'hE0;
            16'd22739: data <= 8'h07;
            16'd22740: data <= 8'hE0;
            16'd22741: data <= 8'h07;
            16'd22742: data <= 8'hE0;
            16'd22743: data <= 8'h07;
            16'd22744: data <= 8'hE0;
            16'd22745: data <= 8'h07;
            16'd22746: data <= 8'hE0;
            16'd22747: data <= 8'h07;
            16'd22748: data <= 8'hE0;
            16'd22749: data <= 8'h07;
            16'd22750: data <= 8'hE0;
            16'd22751: data <= 8'h07;
            16'd22752: data <= 8'hE0;
            16'd22753: data <= 8'h07;
            16'd22754: data <= 8'hE0;
            16'd22755: data <= 8'h07;
            16'd22756: data <= 8'hE0;
            16'd22757: data <= 8'h07;
            16'd22758: data <= 8'hE0;
            16'd22759: data <= 8'h07;
            16'd22760: data <= 8'hFF;
            16'd22761: data <= 8'hFF;
            16'd22762: data <= 8'hE0;
            16'd22763: data <= 8'h07;
            16'd22764: data <= 8'hE0;
            16'd22765: data <= 8'h07;
            16'd22766: data <= 8'hE0;
            16'd22767: data <= 8'h07;
            16'd22768: data <= 8'hE0;
            16'd22769: data <= 8'h07;
            16'd22770: data <= 8'hE0;
            16'd22771: data <= 8'h07;
            16'd22772: data <= 8'hE0;
            16'd22773: data <= 8'h07;
            16'd22774: data <= 8'hE0;
            16'd22775: data <= 8'h07;
            16'd22776: data <= 8'hE0;
            16'd22777: data <= 8'h07;
            16'd22778: data <= 8'hE0;
            16'd22779: data <= 8'h07;
            16'd22780: data <= 8'hE0;
            16'd22781: data <= 8'h07;
            16'd22782: data <= 8'hE0;
            16'd22783: data <= 8'h07;
            16'd22784: data <= 8'hE0;
            16'd22785: data <= 8'h07;
            16'd22786: data <= 8'hE0;
            16'd22787: data <= 8'h07;
            16'd22788: data <= 8'hE0;
            16'd22789: data <= 8'h07;
            16'd22790: data <= 8'hE0;
            16'd22791: data <= 8'h07;
            16'd22792: data <= 8'hE0;
            16'd22793: data <= 8'h07;
            16'd22794: data <= 8'hE0;
            16'd22795: data <= 8'h07;
            16'd22796: data <= 8'hE0;
            16'd22797: data <= 8'h07;
            16'd22798: data <= 8'hE0;
            16'd22799: data <= 8'h07;
            16'd22800: data <= 8'hFF;
            16'd22801: data <= 8'hFF;
            16'd22802: data <= 8'hE0;
            16'd22803: data <= 8'h07;
            16'd22804: data <= 8'hE0;
            16'd22805: data <= 8'h07;
            16'd22806: data <= 8'hE0;
            16'd22807: data <= 8'h07;
            16'd22808: data <= 8'hE0;
            16'd22809: data <= 8'h07;
            16'd22810: data <= 8'hE0;
            16'd22811: data <= 8'h07;
            16'd22812: data <= 8'hE0;
            16'd22813: data <= 8'h07;
            16'd22814: data <= 8'hE0;
            16'd22815: data <= 8'h07;
            16'd22816: data <= 8'hE0;
            16'd22817: data <= 8'h07;
            16'd22818: data <= 8'hE0;
            16'd22819: data <= 8'h07;
            16'd22820: data <= 8'hE0;
            16'd22821: data <= 8'h07;
            16'd22822: data <= 8'hE0;
            16'd22823: data <= 8'h07;
            16'd22824: data <= 8'hE0;
            16'd22825: data <= 8'h07;
            16'd22826: data <= 8'hE0;
            16'd22827: data <= 8'h07;
            16'd22828: data <= 8'hE0;
            16'd22829: data <= 8'h07;
            16'd22830: data <= 8'hE0;
            16'd22831: data <= 8'h07;
            16'd22832: data <= 8'hE0;
            16'd22833: data <= 8'h07;
            16'd22834: data <= 8'hE0;
            16'd22835: data <= 8'h07;
            16'd22836: data <= 8'hE0;
            16'd22837: data <= 8'h07;
            16'd22838: data <= 8'hE0;
            16'd22839: data <= 8'h07;
            16'd22840: data <= 8'hFF;
            16'd22841: data <= 8'hFF;
            16'd22842: data <= 8'hE0;
            16'd22843: data <= 8'h07;
            16'd22844: data <= 8'hE0;
            16'd22845: data <= 8'h07;
            16'd22846: data <= 8'hE0;
            16'd22847: data <= 8'h07;
            16'd22848: data <= 8'hE0;
            16'd22849: data <= 8'h07;
            16'd22850: data <= 8'hE0;
            16'd22851: data <= 8'h07;
            16'd22852: data <= 8'hE0;
            16'd22853: data <= 8'h07;
            16'd22854: data <= 8'hE0;
            16'd22855: data <= 8'h07;
            16'd22856: data <= 8'hE0;
            16'd22857: data <= 8'h07;
            16'd22858: data <= 8'hE0;
            16'd22859: data <= 8'h07;
            16'd22860: data <= 8'hE0;
            16'd22861: data <= 8'h07;
            16'd22862: data <= 8'hE0;
            16'd22863: data <= 8'h07;
            16'd22864: data <= 8'hE0;
            16'd22865: data <= 8'h07;
            16'd22866: data <= 8'hE0;
            16'd22867: data <= 8'h07;
            16'd22868: data <= 8'hE0;
            16'd22869: data <= 8'h07;
            16'd22870: data <= 8'hE0;
            16'd22871: data <= 8'h07;
            16'd22872: data <= 8'hE0;
            16'd22873: data <= 8'h07;
            16'd22874: data <= 8'hE0;
            16'd22875: data <= 8'h07;
            16'd22876: data <= 8'hE0;
            16'd22877: data <= 8'h07;
            16'd22878: data <= 8'hE0;
            16'd22879: data <= 8'h07;
            16'd22880: data <= 8'hFF;
            16'd22881: data <= 8'hFF;
            16'd22882: data <= 8'hE0;
            16'd22883: data <= 8'h07;
            16'd22884: data <= 8'hE0;
            16'd22885: data <= 8'h07;
            16'd22886: data <= 8'hE0;
            16'd22887: data <= 8'h07;
            16'd22888: data <= 8'hE0;
            16'd22889: data <= 8'h07;
            16'd22890: data <= 8'hE0;
            16'd22891: data <= 8'h07;
            16'd22892: data <= 8'hE0;
            16'd22893: data <= 8'h07;
            16'd22894: data <= 8'hE0;
            16'd22895: data <= 8'h07;
            16'd22896: data <= 8'hE0;
            16'd22897: data <= 8'h07;
            16'd22898: data <= 8'hE0;
            16'd22899: data <= 8'h07;
            16'd22900: data <= 8'hE0;
            16'd22901: data <= 8'h07;
            16'd22902: data <= 8'hE0;
            16'd22903: data <= 8'h07;
            16'd22904: data <= 8'hE0;
            16'd22905: data <= 8'h07;
            16'd22906: data <= 8'hE0;
            16'd22907: data <= 8'h07;
            16'd22908: data <= 8'hE0;
            16'd22909: data <= 8'h07;
            16'd22910: data <= 8'hE0;
            16'd22911: data <= 8'h07;
            16'd22912: data <= 8'hE0;
            16'd22913: data <= 8'h07;
            16'd22914: data <= 8'hE0;
            16'd22915: data <= 8'h07;
            16'd22916: data <= 8'hE0;
            16'd22917: data <= 8'h07;
            16'd22918: data <= 8'hE0;
            16'd22919: data <= 8'h07;
            16'd22920: data <= 8'hFF;
            16'd22921: data <= 8'hFF;
            16'd22922: data <= 8'hE0;
            16'd22923: data <= 8'h07;
            16'd22924: data <= 8'hE0;
            16'd22925: data <= 8'h07;
            16'd22926: data <= 8'hE0;
            16'd22927: data <= 8'h07;
            16'd22928: data <= 8'hE0;
            16'd22929: data <= 8'h07;
            16'd22930: data <= 8'hE0;
            16'd22931: data <= 8'h07;
            16'd22932: data <= 8'hE0;
            16'd22933: data <= 8'h07;
            16'd22934: data <= 8'hE0;
            16'd22935: data <= 8'h07;
            16'd22936: data <= 8'hE0;
            16'd22937: data <= 8'h07;
            16'd22938: data <= 8'hE0;
            16'd22939: data <= 8'h07;
            16'd22940: data <= 8'hE0;
            16'd22941: data <= 8'h07;
            16'd22942: data <= 8'hE0;
            16'd22943: data <= 8'h07;
            16'd22944: data <= 8'hE0;
            16'd22945: data <= 8'h07;
            16'd22946: data <= 8'hE0;
            16'd22947: data <= 8'h07;
            16'd22948: data <= 8'hE0;
            16'd22949: data <= 8'h07;
            16'd22950: data <= 8'hE0;
            16'd22951: data <= 8'h07;
            16'd22952: data <= 8'hE0;
            16'd22953: data <= 8'h07;
            16'd22954: data <= 8'hE0;
            16'd22955: data <= 8'h07;
            16'd22956: data <= 8'hE0;
            16'd22957: data <= 8'h07;
            16'd22958: data <= 8'hE0;
            16'd22959: data <= 8'h07;
            16'd22960: data <= 8'hFF;
            16'd22961: data <= 8'hFF;
            16'd22962: data <= 8'hE0;
            16'd22963: data <= 8'h07;
            16'd22964: data <= 8'hE0;
            16'd22965: data <= 8'h07;
            16'd22966: data <= 8'hE0;
            16'd22967: data <= 8'h07;
            16'd22968: data <= 8'hE0;
            16'd22969: data <= 8'h07;
            16'd22970: data <= 8'hE0;
            16'd22971: data <= 8'h07;
            16'd22972: data <= 8'hE0;
            16'd22973: data <= 8'h07;
            16'd22974: data <= 8'hE0;
            16'd22975: data <= 8'h07;
            16'd22976: data <= 8'hE0;
            16'd22977: data <= 8'h07;
            16'd22978: data <= 8'hE0;
            16'd22979: data <= 8'h07;
            16'd22980: data <= 8'hE0;
            16'd22981: data <= 8'h07;
            16'd22982: data <= 8'hE0;
            16'd22983: data <= 8'h07;
            16'd22984: data <= 8'hE0;
            16'd22985: data <= 8'h07;
            16'd22986: data <= 8'hE0;
            16'd22987: data <= 8'h07;
            16'd22988: data <= 8'hE0;
            16'd22989: data <= 8'h07;
            16'd22990: data <= 8'hE0;
            16'd22991: data <= 8'h07;
            16'd22992: data <= 8'hE0;
            16'd22993: data <= 8'h07;
            16'd22994: data <= 8'hE0;
            16'd22995: data <= 8'h07;
            16'd22996: data <= 8'hE0;
            16'd22997: data <= 8'h07;
            16'd22998: data <= 8'hE0;
            16'd22999: data <= 8'h07;
            16'd23000: data <= 8'hFF;
            16'd23001: data <= 8'hFF;
            16'd23002: data <= 8'hE0;
            16'd23003: data <= 8'h07;
            16'd23004: data <= 8'hE0;
            16'd23005: data <= 8'h07;
            16'd23006: data <= 8'hE0;
            16'd23007: data <= 8'h07;
            16'd23008: data <= 8'hE0;
            16'd23009: data <= 8'h07;
            16'd23010: data <= 8'hE0;
            16'd23011: data <= 8'h07;
            16'd23012: data <= 8'hE0;
            16'd23013: data <= 8'h07;
            16'd23014: data <= 8'hE0;
            16'd23015: data <= 8'h07;
            16'd23016: data <= 8'hE0;
            16'd23017: data <= 8'h07;
            16'd23018: data <= 8'hE0;
            16'd23019: data <= 8'h07;
            16'd23020: data <= 8'hE0;
            16'd23021: data <= 8'h07;
            16'd23022: data <= 8'hE0;
            16'd23023: data <= 8'h07;
            16'd23024: data <= 8'hE0;
            16'd23025: data <= 8'h07;
            16'd23026: data <= 8'hE0;
            16'd23027: data <= 8'h07;
            16'd23028: data <= 8'hE0;
            16'd23029: data <= 8'h07;
            16'd23030: data <= 8'hE0;
            16'd23031: data <= 8'h07;
            16'd23032: data <= 8'hE0;
            16'd23033: data <= 8'h07;
            16'd23034: data <= 8'hE0;
            16'd23035: data <= 8'h07;
            16'd23036: data <= 8'hE0;
            16'd23037: data <= 8'h07;
            16'd23038: data <= 8'hE0;
            16'd23039: data <= 8'h07;
            16'd23040: data <= 8'hFF;
            16'd23041: data <= 8'hFF;
            16'd23042: data <= 8'hE0;
            16'd23043: data <= 8'h07;
            16'd23044: data <= 8'hE0;
            16'd23045: data <= 8'h07;
            16'd23046: data <= 8'hE0;
            16'd23047: data <= 8'h07;
            16'd23048: data <= 8'hE0;
            16'd23049: data <= 8'h07;
            16'd23050: data <= 8'hE0;
            16'd23051: data <= 8'h07;
            16'd23052: data <= 8'hE0;
            16'd23053: data <= 8'h07;
            16'd23054: data <= 8'hE0;
            16'd23055: data <= 8'h07;
            16'd23056: data <= 8'hE0;
            16'd23057: data <= 8'h07;
            16'd23058: data <= 8'hE0;
            16'd23059: data <= 8'h07;
            16'd23060: data <= 8'hE0;
            16'd23061: data <= 8'h07;
            16'd23062: data <= 8'hE0;
            16'd23063: data <= 8'h07;
            16'd23064: data <= 8'hE0;
            16'd23065: data <= 8'h07;
            16'd23066: data <= 8'hE0;
            16'd23067: data <= 8'h07;
            16'd23068: data <= 8'hE0;
            16'd23069: data <= 8'h07;
            16'd23070: data <= 8'hE0;
            16'd23071: data <= 8'h07;
            16'd23072: data <= 8'hE0;
            16'd23073: data <= 8'h07;
            16'd23074: data <= 8'hE0;
            16'd23075: data <= 8'h07;
            16'd23076: data <= 8'hE0;
            16'd23077: data <= 8'h07;
            16'd23078: data <= 8'hE0;
            16'd23079: data <= 8'h07;
            16'd23080: data <= 8'hFF;
            16'd23081: data <= 8'hFF;
            16'd23082: data <= 8'hE0;
            16'd23083: data <= 8'h07;
            16'd23084: data <= 8'hE0;
            16'd23085: data <= 8'h07;
            16'd23086: data <= 8'hE0;
            16'd23087: data <= 8'h07;
            16'd23088: data <= 8'hE0;
            16'd23089: data <= 8'h07;
            16'd23090: data <= 8'hE0;
            16'd23091: data <= 8'h07;
            16'd23092: data <= 8'hE0;
            16'd23093: data <= 8'h07;
            16'd23094: data <= 8'hE0;
            16'd23095: data <= 8'h07;
            16'd23096: data <= 8'hE0;
            16'd23097: data <= 8'h07;
            16'd23098: data <= 8'hE0;
            16'd23099: data <= 8'h07;
            16'd23100: data <= 8'hE0;
            16'd23101: data <= 8'h07;
            16'd23102: data <= 8'hE0;
            16'd23103: data <= 8'h07;
            16'd23104: data <= 8'hE0;
            16'd23105: data <= 8'h07;
            16'd23106: data <= 8'hE0;
            16'd23107: data <= 8'h07;
            16'd23108: data <= 8'hE0;
            16'd23109: data <= 8'h07;
            16'd23110: data <= 8'hE0;
            16'd23111: data <= 8'h07;
            16'd23112: data <= 8'hE0;
            16'd23113: data <= 8'h07;
            16'd23114: data <= 8'hE0;
            16'd23115: data <= 8'h07;
            16'd23116: data <= 8'hE0;
            16'd23117: data <= 8'h07;
            16'd23118: data <= 8'hE0;
            16'd23119: data <= 8'h07;
            16'd23120: data <= 8'hFF;
            16'd23121: data <= 8'hFF;
            16'd23122: data <= 8'hE0;
            16'd23123: data <= 8'h07;
            16'd23124: data <= 8'hE0;
            16'd23125: data <= 8'h07;
            16'd23126: data <= 8'hE0;
            16'd23127: data <= 8'h07;
            16'd23128: data <= 8'hE0;
            16'd23129: data <= 8'h07;
            16'd23130: data <= 8'hE0;
            16'd23131: data <= 8'h07;
            16'd23132: data <= 8'hE0;
            16'd23133: data <= 8'h07;
            16'd23134: data <= 8'hE0;
            16'd23135: data <= 8'h07;
            16'd23136: data <= 8'hE0;
            16'd23137: data <= 8'h07;
            16'd23138: data <= 8'hE0;
            16'd23139: data <= 8'h07;
            16'd23140: data <= 8'hE0;
            16'd23141: data <= 8'h07;
            16'd23142: data <= 8'hE0;
            16'd23143: data <= 8'h07;
            16'd23144: data <= 8'hE0;
            16'd23145: data <= 8'h07;
            16'd23146: data <= 8'hE0;
            16'd23147: data <= 8'h07;
            16'd23148: data <= 8'hE0;
            16'd23149: data <= 8'h07;
            16'd23150: data <= 8'hE0;
            16'd23151: data <= 8'h07;
            16'd23152: data <= 8'hE0;
            16'd23153: data <= 8'h07;
            16'd23154: data <= 8'hE0;
            16'd23155: data <= 8'h07;
            16'd23156: data <= 8'hE0;
            16'd23157: data <= 8'h07;
            16'd23158: data <= 8'hE0;
            16'd23159: data <= 8'h07;
            16'd23160: data <= 8'hFF;
            16'd23161: data <= 8'hFF;
            16'd23162: data <= 8'hE0;
            16'd23163: data <= 8'h07;
            16'd23164: data <= 8'hE0;
            16'd23165: data <= 8'h07;
            16'd23166: data <= 8'hE0;
            16'd23167: data <= 8'h07;
            16'd23168: data <= 8'hE0;
            16'd23169: data <= 8'h07;
            16'd23170: data <= 8'hE0;
            16'd23171: data <= 8'h07;
            16'd23172: data <= 8'hE0;
            16'd23173: data <= 8'h07;
            16'd23174: data <= 8'hE0;
            16'd23175: data <= 8'h07;
            16'd23176: data <= 8'hE0;
            16'd23177: data <= 8'h07;
            16'd23178: data <= 8'hE0;
            16'd23179: data <= 8'h07;
            16'd23180: data <= 8'hE0;
            16'd23181: data <= 8'h07;
            16'd23182: data <= 8'hE0;
            16'd23183: data <= 8'h07;
            16'd23184: data <= 8'hE0;
            16'd23185: data <= 8'h07;
            16'd23186: data <= 8'hE0;
            16'd23187: data <= 8'h07;
            16'd23188: data <= 8'hE0;
            16'd23189: data <= 8'h07;
            16'd23190: data <= 8'hE0;
            16'd23191: data <= 8'h07;
            16'd23192: data <= 8'hE0;
            16'd23193: data <= 8'h07;
            16'd23194: data <= 8'hE0;
            16'd23195: data <= 8'h07;
            16'd23196: data <= 8'hE0;
            16'd23197: data <= 8'h07;
            16'd23198: data <= 8'hE0;
            16'd23199: data <= 8'h07;
            16'd23200: data <= 8'hFF;
            16'd23201: data <= 8'hFF;
            16'd23202: data <= 8'hE0;
            16'd23203: data <= 8'h07;
            16'd23204: data <= 8'hE0;
            16'd23205: data <= 8'h07;
            16'd23206: data <= 8'hE0;
            16'd23207: data <= 8'h07;
            16'd23208: data <= 8'hE0;
            16'd23209: data <= 8'h07;
            16'd23210: data <= 8'hE0;
            16'd23211: data <= 8'h07;
            16'd23212: data <= 8'hE0;
            16'd23213: data <= 8'h07;
            16'd23214: data <= 8'hE0;
            16'd23215: data <= 8'h07;
            16'd23216: data <= 8'hE0;
            16'd23217: data <= 8'h07;
            16'd23218: data <= 8'hE0;
            16'd23219: data <= 8'h07;
            16'd23220: data <= 8'hE0;
            16'd23221: data <= 8'h07;
            16'd23222: data <= 8'hE0;
            16'd23223: data <= 8'h07;
            16'd23224: data <= 8'hE0;
            16'd23225: data <= 8'h07;
            16'd23226: data <= 8'hE0;
            16'd23227: data <= 8'h07;
            16'd23228: data <= 8'hE0;
            16'd23229: data <= 8'h07;
            16'd23230: data <= 8'hE0;
            16'd23231: data <= 8'h07;
            16'd23232: data <= 8'hE0;
            16'd23233: data <= 8'h07;
            16'd23234: data <= 8'hE0;
            16'd23235: data <= 8'h07;
            16'd23236: data <= 8'hE0;
            16'd23237: data <= 8'h07;
            16'd23238: data <= 8'hE0;
            16'd23239: data <= 8'h07;
            16'd23240: data <= 8'hFF;
            16'd23241: data <= 8'hFF;
            16'd23242: data <= 8'hE0;
            16'd23243: data <= 8'h07;
            16'd23244: data <= 8'hE0;
            16'd23245: data <= 8'h07;
            16'd23246: data <= 8'hE0;
            16'd23247: data <= 8'h07;
            16'd23248: data <= 8'hE0;
            16'd23249: data <= 8'h07;
            16'd23250: data <= 8'hE0;
            16'd23251: data <= 8'h07;
            16'd23252: data <= 8'hE0;
            16'd23253: data <= 8'h07;
            16'd23254: data <= 8'hE0;
            16'd23255: data <= 8'h07;
            16'd23256: data <= 8'hE0;
            16'd23257: data <= 8'h07;
            16'd23258: data <= 8'hE0;
            16'd23259: data <= 8'h07;
            16'd23260: data <= 8'hE0;
            16'd23261: data <= 8'h07;
            16'd23262: data <= 8'hE0;
            16'd23263: data <= 8'h07;
            16'd23264: data <= 8'hE0;
            16'd23265: data <= 8'h07;
            16'd23266: data <= 8'hE0;
            16'd23267: data <= 8'h07;
            16'd23268: data <= 8'hE0;
            16'd23269: data <= 8'h07;
            16'd23270: data <= 8'hE0;
            16'd23271: data <= 8'h07;
            16'd23272: data <= 8'hE0;
            16'd23273: data <= 8'h07;
            16'd23274: data <= 8'hE0;
            16'd23275: data <= 8'h07;
            16'd23276: data <= 8'hE0;
            16'd23277: data <= 8'h07;
            16'd23278: data <= 8'hE0;
            16'd23279: data <= 8'h07;
            16'd23280: data <= 8'hFF;
            16'd23281: data <= 8'hFF;
            16'd23282: data <= 8'hE0;
            16'd23283: data <= 8'h07;
            16'd23284: data <= 8'hE0;
            16'd23285: data <= 8'h07;
            16'd23286: data <= 8'hE0;
            16'd23287: data <= 8'h07;
            16'd23288: data <= 8'hE0;
            16'd23289: data <= 8'h07;
            16'd23290: data <= 8'hE0;
            16'd23291: data <= 8'h07;
            16'd23292: data <= 8'hE0;
            16'd23293: data <= 8'h07;
            16'd23294: data <= 8'hE0;
            16'd23295: data <= 8'h07;
            16'd23296: data <= 8'hE0;
            16'd23297: data <= 8'h07;
            16'd23298: data <= 8'hE0;
            16'd23299: data <= 8'h07;
            16'd23300: data <= 8'hE0;
            16'd23301: data <= 8'h07;
            16'd23302: data <= 8'hE0;
            16'd23303: data <= 8'h07;
            16'd23304: data <= 8'hE0;
            16'd23305: data <= 8'h07;
            16'd23306: data <= 8'hE0;
            16'd23307: data <= 8'h07;
            16'd23308: data <= 8'hE0;
            16'd23309: data <= 8'h07;
            16'd23310: data <= 8'hE0;
            16'd23311: data <= 8'h07;
            16'd23312: data <= 8'hE0;
            16'd23313: data <= 8'h07;
            16'd23314: data <= 8'hE0;
            16'd23315: data <= 8'h07;
            16'd23316: data <= 8'hE0;
            16'd23317: data <= 8'h07;
            16'd23318: data <= 8'hE0;
            16'd23319: data <= 8'h07;
            16'd23320: data <= 8'hFF;
            16'd23321: data <= 8'hFF;
            16'd23322: data <= 8'hE0;
            16'd23323: data <= 8'h07;
            16'd23324: data <= 8'hE0;
            16'd23325: data <= 8'h07;
            16'd23326: data <= 8'hE0;
            16'd23327: data <= 8'h07;
            16'd23328: data <= 8'hE0;
            16'd23329: data <= 8'h07;
            16'd23330: data <= 8'hE0;
            16'd23331: data <= 8'h07;
            16'd23332: data <= 8'hE0;
            16'd23333: data <= 8'h07;
            16'd23334: data <= 8'hE0;
            16'd23335: data <= 8'h07;
            16'd23336: data <= 8'hE0;
            16'd23337: data <= 8'h07;
            16'd23338: data <= 8'hE0;
            16'd23339: data <= 8'h07;
            16'd23340: data <= 8'hE0;
            16'd23341: data <= 8'h07;
            16'd23342: data <= 8'hE0;
            16'd23343: data <= 8'h07;
            16'd23344: data <= 8'hE0;
            16'd23345: data <= 8'h07;
            16'd23346: data <= 8'hE0;
            16'd23347: data <= 8'h07;
            16'd23348: data <= 8'hE0;
            16'd23349: data <= 8'h07;
            16'd23350: data <= 8'hE0;
            16'd23351: data <= 8'h07;
            16'd23352: data <= 8'hE0;
            16'd23353: data <= 8'h07;
            16'd23354: data <= 8'hE0;
            16'd23355: data <= 8'h07;
            16'd23356: data <= 8'hE0;
            16'd23357: data <= 8'h07;
            16'd23358: data <= 8'hE0;
            16'd23359: data <= 8'h07;
            16'd23360: data <= 8'hFF;
            16'd23361: data <= 8'hFF;
            16'd23362: data <= 8'hE0;
            16'd23363: data <= 8'h07;
            16'd23364: data <= 8'hE0;
            16'd23365: data <= 8'h07;
            16'd23366: data <= 8'hE0;
            16'd23367: data <= 8'h07;
            16'd23368: data <= 8'hE0;
            16'd23369: data <= 8'h07;
            16'd23370: data <= 8'hE0;
            16'd23371: data <= 8'h07;
            16'd23372: data <= 8'hE0;
            16'd23373: data <= 8'h07;
            16'd23374: data <= 8'hE0;
            16'd23375: data <= 8'h07;
            16'd23376: data <= 8'hE0;
            16'd23377: data <= 8'h07;
            16'd23378: data <= 8'hE0;
            16'd23379: data <= 8'h07;
            16'd23380: data <= 8'hE0;
            16'd23381: data <= 8'h07;
            16'd23382: data <= 8'hE0;
            16'd23383: data <= 8'h07;
            16'd23384: data <= 8'hE0;
            16'd23385: data <= 8'h07;
            16'd23386: data <= 8'hE0;
            16'd23387: data <= 8'h07;
            16'd23388: data <= 8'hE0;
            16'd23389: data <= 8'h07;
            16'd23390: data <= 8'hE0;
            16'd23391: data <= 8'h07;
            16'd23392: data <= 8'hE0;
            16'd23393: data <= 8'h07;
            16'd23394: data <= 8'hE0;
            16'd23395: data <= 8'h07;
            16'd23396: data <= 8'hE0;
            16'd23397: data <= 8'h07;
            16'd23398: data <= 8'hE0;
            16'd23399: data <= 8'h07;
            16'd23400: data <= 8'hFF;
            16'd23401: data <= 8'hFF;
            16'd23402: data <= 8'hE0;
            16'd23403: data <= 8'h07;
            16'd23404: data <= 8'hE0;
            16'd23405: data <= 8'h07;
            16'd23406: data <= 8'hE0;
            16'd23407: data <= 8'h07;
            16'd23408: data <= 8'hE0;
            16'd23409: data <= 8'h07;
            16'd23410: data <= 8'hE0;
            16'd23411: data <= 8'h07;
            16'd23412: data <= 8'hE0;
            16'd23413: data <= 8'h07;
            16'd23414: data <= 8'hE0;
            16'd23415: data <= 8'h07;
            16'd23416: data <= 8'hE0;
            16'd23417: data <= 8'h07;
            16'd23418: data <= 8'hE0;
            16'd23419: data <= 8'h07;
            16'd23420: data <= 8'hE0;
            16'd23421: data <= 8'h07;
            16'd23422: data <= 8'hE0;
            16'd23423: data <= 8'h07;
            16'd23424: data <= 8'hE0;
            16'd23425: data <= 8'h07;
            16'd23426: data <= 8'hE0;
            16'd23427: data <= 8'h07;
            16'd23428: data <= 8'hE0;
            16'd23429: data <= 8'h07;
            16'd23430: data <= 8'hE0;
            16'd23431: data <= 8'h07;
            16'd23432: data <= 8'hE0;
            16'd23433: data <= 8'h07;
            16'd23434: data <= 8'hE0;
            16'd23435: data <= 8'h07;
            16'd23436: data <= 8'hE0;
            16'd23437: data <= 8'h07;
            16'd23438: data <= 8'hE0;
            16'd23439: data <= 8'h07;
            16'd23440: data <= 8'hFF;
            16'd23441: data <= 8'hFF;
            16'd23442: data <= 8'hE0;
            16'd23443: data <= 8'h07;
            16'd23444: data <= 8'hE0;
            16'd23445: data <= 8'h07;
            16'd23446: data <= 8'hE0;
            16'd23447: data <= 8'h07;
            16'd23448: data <= 8'hE0;
            16'd23449: data <= 8'h07;
            16'd23450: data <= 8'hE0;
            16'd23451: data <= 8'h07;
            16'd23452: data <= 8'hE0;
            16'd23453: data <= 8'h07;
            16'd23454: data <= 8'hE0;
            16'd23455: data <= 8'h07;
            16'd23456: data <= 8'hE0;
            16'd23457: data <= 8'h07;
            16'd23458: data <= 8'hE0;
            16'd23459: data <= 8'h07;
            16'd23460: data <= 8'hE0;
            16'd23461: data <= 8'h07;
            16'd23462: data <= 8'hE0;
            16'd23463: data <= 8'h07;
            16'd23464: data <= 8'hE0;
            16'd23465: data <= 8'h07;
            16'd23466: data <= 8'hE0;
            16'd23467: data <= 8'h07;
            16'd23468: data <= 8'hE0;
            16'd23469: data <= 8'h07;
            16'd23470: data <= 8'hE0;
            16'd23471: data <= 8'h07;
            16'd23472: data <= 8'hE0;
            16'd23473: data <= 8'h07;
            16'd23474: data <= 8'hE0;
            16'd23475: data <= 8'h07;
            16'd23476: data <= 8'hE0;
            16'd23477: data <= 8'h07;
            16'd23478: data <= 8'hE0;
            16'd23479: data <= 8'h07;
            16'd23480: data <= 8'hFF;
            16'd23481: data <= 8'hFF;
            16'd23482: data <= 8'hE0;
            16'd23483: data <= 8'h07;
            16'd23484: data <= 8'hE0;
            16'd23485: data <= 8'h07;
            16'd23486: data <= 8'hE0;
            16'd23487: data <= 8'h07;
            16'd23488: data <= 8'hE0;
            16'd23489: data <= 8'h07;
            16'd23490: data <= 8'hE0;
            16'd23491: data <= 8'h07;
            16'd23492: data <= 8'hE0;
            16'd23493: data <= 8'h07;
            16'd23494: data <= 8'hE0;
            16'd23495: data <= 8'h07;
            16'd23496: data <= 8'hE0;
            16'd23497: data <= 8'h07;
            16'd23498: data <= 8'hE0;
            16'd23499: data <= 8'h07;
            16'd23500: data <= 8'hE0;
            16'd23501: data <= 8'h07;
            16'd23502: data <= 8'hE0;
            16'd23503: data <= 8'h07;
            16'd23504: data <= 8'hE0;
            16'd23505: data <= 8'h07;
            16'd23506: data <= 8'hE0;
            16'd23507: data <= 8'h07;
            16'd23508: data <= 8'hE0;
            16'd23509: data <= 8'h07;
            16'd23510: data <= 8'hE0;
            16'd23511: data <= 8'h07;
            16'd23512: data <= 8'hE0;
            16'd23513: data <= 8'h07;
            16'd23514: data <= 8'hE0;
            16'd23515: data <= 8'h07;
            16'd23516: data <= 8'hE0;
            16'd23517: data <= 8'h07;
            16'd23518: data <= 8'hE0;
            16'd23519: data <= 8'h07;
            16'd23520: data <= 8'hFF;
            16'd23521: data <= 8'hFF;
            16'd23522: data <= 8'hE0;
            16'd23523: data <= 8'h07;
            16'd23524: data <= 8'hE0;
            16'd23525: data <= 8'h07;
            16'd23526: data <= 8'hE0;
            16'd23527: data <= 8'h07;
            16'd23528: data <= 8'hE0;
            16'd23529: data <= 8'h07;
            16'd23530: data <= 8'hE0;
            16'd23531: data <= 8'h07;
            16'd23532: data <= 8'hE0;
            16'd23533: data <= 8'h07;
            16'd23534: data <= 8'hE0;
            16'd23535: data <= 8'h07;
            16'd23536: data <= 8'hE0;
            16'd23537: data <= 8'h07;
            16'd23538: data <= 8'hE0;
            16'd23539: data <= 8'h07;
            16'd23540: data <= 8'hE0;
            16'd23541: data <= 8'h07;
            16'd23542: data <= 8'hE0;
            16'd23543: data <= 8'h07;
            16'd23544: data <= 8'hE0;
            16'd23545: data <= 8'h07;
            16'd23546: data <= 8'hE0;
            16'd23547: data <= 8'h07;
            16'd23548: data <= 8'hE0;
            16'd23549: data <= 8'h07;
            16'd23550: data <= 8'hE0;
            16'd23551: data <= 8'h07;
            16'd23552: data <= 8'hE0;
            16'd23553: data <= 8'h07;
            16'd23554: data <= 8'hE0;
            16'd23555: data <= 8'h07;
            16'd23556: data <= 8'hE0;
            16'd23557: data <= 8'h07;
            16'd23558: data <= 8'hE0;
            16'd23559: data <= 8'h07;
            16'd23560: data <= 8'hFF;
            16'd23561: data <= 8'hFF;
            16'd23562: data <= 8'hE0;
            16'd23563: data <= 8'h07;
            16'd23564: data <= 8'hE0;
            16'd23565: data <= 8'h07;
            16'd23566: data <= 8'hE0;
            16'd23567: data <= 8'h07;
            16'd23568: data <= 8'hE0;
            16'd23569: data <= 8'h07;
            16'd23570: data <= 8'hE0;
            16'd23571: data <= 8'h07;
            16'd23572: data <= 8'hE0;
            16'd23573: data <= 8'h07;
            16'd23574: data <= 8'hE0;
            16'd23575: data <= 8'h07;
            16'd23576: data <= 8'hE0;
            16'd23577: data <= 8'h07;
            16'd23578: data <= 8'hE0;
            16'd23579: data <= 8'h07;
            16'd23580: data <= 8'hE0;
            16'd23581: data <= 8'h07;
            16'd23582: data <= 8'hE0;
            16'd23583: data <= 8'h07;
            16'd23584: data <= 8'hE0;
            16'd23585: data <= 8'h07;
            16'd23586: data <= 8'hE0;
            16'd23587: data <= 8'h07;
            16'd23588: data <= 8'hE0;
            16'd23589: data <= 8'h07;
            16'd23590: data <= 8'hE0;
            16'd23591: data <= 8'h07;
            16'd23592: data <= 8'hE0;
            16'd23593: data <= 8'h07;
            16'd23594: data <= 8'hE0;
            16'd23595: data <= 8'h07;
            16'd23596: data <= 8'hE0;
            16'd23597: data <= 8'h07;
            16'd23598: data <= 8'hE0;
            16'd23599: data <= 8'h07;
            16'd23600: data <= 8'hFF;
            16'd23601: data <= 8'hFF;
            16'd23602: data <= 8'hE0;
            16'd23603: data <= 8'h07;
            16'd23604: data <= 8'hE0;
            16'd23605: data <= 8'h07;
            16'd23606: data <= 8'hE0;
            16'd23607: data <= 8'h07;
            16'd23608: data <= 8'hE0;
            16'd23609: data <= 8'h07;
            16'd23610: data <= 8'hE0;
            16'd23611: data <= 8'h07;
            16'd23612: data <= 8'hE0;
            16'd23613: data <= 8'h07;
            16'd23614: data <= 8'hE0;
            16'd23615: data <= 8'h07;
            16'd23616: data <= 8'hE0;
            16'd23617: data <= 8'h07;
            16'd23618: data <= 8'hE0;
            16'd23619: data <= 8'h07;
            16'd23620: data <= 8'hE0;
            16'd23621: data <= 8'h07;
            16'd23622: data <= 8'hE0;
            16'd23623: data <= 8'h07;
            16'd23624: data <= 8'hE0;
            16'd23625: data <= 8'h07;
            16'd23626: data <= 8'hE0;
            16'd23627: data <= 8'h07;
            16'd23628: data <= 8'hE0;
            16'd23629: data <= 8'h07;
            16'd23630: data <= 8'hE0;
            16'd23631: data <= 8'h07;
            16'd23632: data <= 8'hE0;
            16'd23633: data <= 8'h07;
            16'd23634: data <= 8'hE0;
            16'd23635: data <= 8'h07;
            16'd23636: data <= 8'hE0;
            16'd23637: data <= 8'h07;
            16'd23638: data <= 8'hE0;
            16'd23639: data <= 8'h07;
            16'd23640: data <= 8'hFF;
            16'd23641: data <= 8'hFF;
            16'd23642: data <= 8'hE0;
            16'd23643: data <= 8'h07;
            16'd23644: data <= 8'hE0;
            16'd23645: data <= 8'h07;
            16'd23646: data <= 8'hE0;
            16'd23647: data <= 8'h07;
            16'd23648: data <= 8'hE0;
            16'd23649: data <= 8'h07;
            16'd23650: data <= 8'hE0;
            16'd23651: data <= 8'h07;
            16'd23652: data <= 8'hE0;
            16'd23653: data <= 8'h07;
            16'd23654: data <= 8'hE0;
            16'd23655: data <= 8'h07;
            16'd23656: data <= 8'hE0;
            16'd23657: data <= 8'h07;
            16'd23658: data <= 8'hE0;
            16'd23659: data <= 8'h07;
            16'd23660: data <= 8'hE0;
            16'd23661: data <= 8'h07;
            16'd23662: data <= 8'hE0;
            16'd23663: data <= 8'h07;
            16'd23664: data <= 8'hE0;
            16'd23665: data <= 8'h07;
            16'd23666: data <= 8'hE0;
            16'd23667: data <= 8'h07;
            16'd23668: data <= 8'hE0;
            16'd23669: data <= 8'h07;
            16'd23670: data <= 8'hE0;
            16'd23671: data <= 8'h07;
            16'd23672: data <= 8'hE0;
            16'd23673: data <= 8'h07;
            16'd23674: data <= 8'hE0;
            16'd23675: data <= 8'h07;
            16'd23676: data <= 8'hE0;
            16'd23677: data <= 8'h07;
            16'd23678: data <= 8'hE0;
            16'd23679: data <= 8'h07;
            16'd23680: data <= 8'hFF;
            16'd23681: data <= 8'hFF;
            16'd23682: data <= 8'hE0;
            16'd23683: data <= 8'h07;
            16'd23684: data <= 8'hE0;
            16'd23685: data <= 8'h07;
            16'd23686: data <= 8'hE0;
            16'd23687: data <= 8'h07;
            16'd23688: data <= 8'hE0;
            16'd23689: data <= 8'h07;
            16'd23690: data <= 8'hE0;
            16'd23691: data <= 8'h07;
            16'd23692: data <= 8'hE0;
            16'd23693: data <= 8'h07;
            16'd23694: data <= 8'hE0;
            16'd23695: data <= 8'h07;
            16'd23696: data <= 8'hE0;
            16'd23697: data <= 8'h07;
            16'd23698: data <= 8'hE0;
            16'd23699: data <= 8'h07;
            16'd23700: data <= 8'hE0;
            16'd23701: data <= 8'h07;
            16'd23702: data <= 8'hE0;
            16'd23703: data <= 8'h07;
            16'd23704: data <= 8'hE0;
            16'd23705: data <= 8'h07;
            16'd23706: data <= 8'hE0;
            16'd23707: data <= 8'h07;
            16'd23708: data <= 8'hE0;
            16'd23709: data <= 8'h07;
            16'd23710: data <= 8'hE0;
            16'd23711: data <= 8'h07;
            16'd23712: data <= 8'hE0;
            16'd23713: data <= 8'h07;
            16'd23714: data <= 8'hE0;
            16'd23715: data <= 8'h07;
            16'd23716: data <= 8'hE0;
            16'd23717: data <= 8'h07;
            16'd23718: data <= 8'hE0;
            16'd23719: data <= 8'h07;
            16'd23720: data <= 8'hFF;
            16'd23721: data <= 8'hFF;
            16'd23722: data <= 8'hE0;
            16'd23723: data <= 8'h07;
            16'd23724: data <= 8'hE0;
            16'd23725: data <= 8'h07;
            16'd23726: data <= 8'hE0;
            16'd23727: data <= 8'h07;
            16'd23728: data <= 8'hE0;
            16'd23729: data <= 8'h07;
            16'd23730: data <= 8'hE0;
            16'd23731: data <= 8'h07;
            16'd23732: data <= 8'hE0;
            16'd23733: data <= 8'h07;
            16'd23734: data <= 8'hE0;
            16'd23735: data <= 8'h07;
            16'd23736: data <= 8'hE0;
            16'd23737: data <= 8'h07;
            16'd23738: data <= 8'hE0;
            16'd23739: data <= 8'h07;
            16'd23740: data <= 8'hE0;
            16'd23741: data <= 8'h07;
            16'd23742: data <= 8'hE0;
            16'd23743: data <= 8'h07;
            16'd23744: data <= 8'hE0;
            16'd23745: data <= 8'h07;
            16'd23746: data <= 8'hE0;
            16'd23747: data <= 8'h07;
            16'd23748: data <= 8'hE0;
            16'd23749: data <= 8'h07;
            16'd23750: data <= 8'hE0;
            16'd23751: data <= 8'h07;
            16'd23752: data <= 8'hE0;
            16'd23753: data <= 8'h07;
            16'd23754: data <= 8'hE0;
            16'd23755: data <= 8'h07;
            16'd23756: data <= 8'hE0;
            16'd23757: data <= 8'h07;
            16'd23758: data <= 8'hE0;
            16'd23759: data <= 8'h07;
            16'd23760: data <= 8'hFF;
            16'd23761: data <= 8'hFF;
            16'd23762: data <= 8'hE0;
            16'd23763: data <= 8'h07;
            16'd23764: data <= 8'hE0;
            16'd23765: data <= 8'h07;
            16'd23766: data <= 8'hE0;
            16'd23767: data <= 8'h07;
            16'd23768: data <= 8'hE0;
            16'd23769: data <= 8'h07;
            16'd23770: data <= 8'hE0;
            16'd23771: data <= 8'h07;
            16'd23772: data <= 8'hE0;
            16'd23773: data <= 8'h07;
            16'd23774: data <= 8'hE0;
            16'd23775: data <= 8'h07;
            16'd23776: data <= 8'hE0;
            16'd23777: data <= 8'h07;
            16'd23778: data <= 8'hE0;
            16'd23779: data <= 8'h07;
            16'd23780: data <= 8'hE0;
            16'd23781: data <= 8'h07;
            16'd23782: data <= 8'hE0;
            16'd23783: data <= 8'h07;
            16'd23784: data <= 8'hE0;
            16'd23785: data <= 8'h07;
            16'd23786: data <= 8'hE0;
            16'd23787: data <= 8'h07;
            16'd23788: data <= 8'hE0;
            16'd23789: data <= 8'h07;
            16'd23790: data <= 8'hE0;
            16'd23791: data <= 8'h07;
            16'd23792: data <= 8'hE0;
            16'd23793: data <= 8'h07;
            16'd23794: data <= 8'hE0;
            16'd23795: data <= 8'h07;
            16'd23796: data <= 8'hE0;
            16'd23797: data <= 8'h07;
            16'd23798: data <= 8'hE0;
            16'd23799: data <= 8'h07;
            16'd23800: data <= 8'hFF;
            16'd23801: data <= 8'hFF;
            16'd23802: data <= 8'hE0;
            16'd23803: data <= 8'h07;
            16'd23804: data <= 8'hE0;
            16'd23805: data <= 8'h07;
            16'd23806: data <= 8'hE0;
            16'd23807: data <= 8'h07;
            16'd23808: data <= 8'hE0;
            16'd23809: data <= 8'h07;
            16'd23810: data <= 8'hE0;
            16'd23811: data <= 8'h07;
            16'd23812: data <= 8'hE0;
            16'd23813: data <= 8'h07;
            16'd23814: data <= 8'hE0;
            16'd23815: data <= 8'h07;
            16'd23816: data <= 8'hE0;
            16'd23817: data <= 8'h07;
            16'd23818: data <= 8'hE0;
            16'd23819: data <= 8'h07;
            16'd23820: data <= 8'hE0;
            16'd23821: data <= 8'h07;
            16'd23822: data <= 8'hE0;
            16'd23823: data <= 8'h07;
            16'd23824: data <= 8'hE0;
            16'd23825: data <= 8'h07;
            16'd23826: data <= 8'hE0;
            16'd23827: data <= 8'h07;
            16'd23828: data <= 8'hE0;
            16'd23829: data <= 8'h07;
            16'd23830: data <= 8'hE0;
            16'd23831: data <= 8'h07;
            16'd23832: data <= 8'hE0;
            16'd23833: data <= 8'h07;
            16'd23834: data <= 8'hE0;
            16'd23835: data <= 8'h07;
            16'd23836: data <= 8'hE0;
            16'd23837: data <= 8'h07;
            16'd23838: data <= 8'hE0;
            16'd23839: data <= 8'h07;
            16'd23840: data <= 8'hFF;
            16'd23841: data <= 8'hFF;
            16'd23842: data <= 8'hE0;
            16'd23843: data <= 8'h07;
            16'd23844: data <= 8'hE0;
            16'd23845: data <= 8'h07;
            16'd23846: data <= 8'hE0;
            16'd23847: data <= 8'h07;
            16'd23848: data <= 8'hE0;
            16'd23849: data <= 8'h07;
            16'd23850: data <= 8'hE0;
            16'd23851: data <= 8'h07;
            16'd23852: data <= 8'hE0;
            16'd23853: data <= 8'h07;
            16'd23854: data <= 8'hE0;
            16'd23855: data <= 8'h07;
            16'd23856: data <= 8'hE0;
            16'd23857: data <= 8'h07;
            16'd23858: data <= 8'hE0;
            16'd23859: data <= 8'h07;
            16'd23860: data <= 8'hE0;
            16'd23861: data <= 8'h07;
            16'd23862: data <= 8'hE0;
            16'd23863: data <= 8'h07;
            16'd23864: data <= 8'hE0;
            16'd23865: data <= 8'h07;
            16'd23866: data <= 8'hE0;
            16'd23867: data <= 8'h07;
            16'd23868: data <= 8'hE0;
            16'd23869: data <= 8'h07;
            16'd23870: data <= 8'hE0;
            16'd23871: data <= 8'h07;
            16'd23872: data <= 8'hE0;
            16'd23873: data <= 8'h07;
            16'd23874: data <= 8'hE0;
            16'd23875: data <= 8'h07;
            16'd23876: data <= 8'hE0;
            16'd23877: data <= 8'h07;
            16'd23878: data <= 8'hE0;
            16'd23879: data <= 8'h07;
            16'd23880: data <= 8'hFF;
            16'd23881: data <= 8'hFF;
            16'd23882: data <= 8'hE0;
            16'd23883: data <= 8'h07;
            16'd23884: data <= 8'hE0;
            16'd23885: data <= 8'h07;
            16'd23886: data <= 8'hE0;
            16'd23887: data <= 8'h07;
            16'd23888: data <= 8'hE0;
            16'd23889: data <= 8'h07;
            16'd23890: data <= 8'hE0;
            16'd23891: data <= 8'h07;
            16'd23892: data <= 8'hE0;
            16'd23893: data <= 8'h07;
            16'd23894: data <= 8'hE0;
            16'd23895: data <= 8'h07;
            16'd23896: data <= 8'hE0;
            16'd23897: data <= 8'h07;
            16'd23898: data <= 8'hE0;
            16'd23899: data <= 8'h07;
            16'd23900: data <= 8'hE0;
            16'd23901: data <= 8'h07;
            16'd23902: data <= 8'hE0;
            16'd23903: data <= 8'h07;
            16'd23904: data <= 8'hE0;
            16'd23905: data <= 8'h07;
            16'd23906: data <= 8'hE0;
            16'd23907: data <= 8'h07;
            16'd23908: data <= 8'hE0;
            16'd23909: data <= 8'h07;
            16'd23910: data <= 8'hE0;
            16'd23911: data <= 8'h07;
            16'd23912: data <= 8'hE0;
            16'd23913: data <= 8'h07;
            16'd23914: data <= 8'hE0;
            16'd23915: data <= 8'h07;
            16'd23916: data <= 8'hE0;
            16'd23917: data <= 8'h07;
            16'd23918: data <= 8'hE0;
            16'd23919: data <= 8'h07;
            16'd23920: data <= 8'hFF;
            16'd23921: data <= 8'hFF;
            16'd23922: data <= 8'hE0;
            16'd23923: data <= 8'h07;
            16'd23924: data <= 8'hE0;
            16'd23925: data <= 8'h07;
            16'd23926: data <= 8'hE0;
            16'd23927: data <= 8'h07;
            16'd23928: data <= 8'hE0;
            16'd23929: data <= 8'h07;
            16'd23930: data <= 8'hE0;
            16'd23931: data <= 8'h07;
            16'd23932: data <= 8'hE0;
            16'd23933: data <= 8'h07;
            16'd23934: data <= 8'hE0;
            16'd23935: data <= 8'h07;
            16'd23936: data <= 8'hE0;
            16'd23937: data <= 8'h07;
            16'd23938: data <= 8'hE0;
            16'd23939: data <= 8'h07;
            16'd23940: data <= 8'hE0;
            16'd23941: data <= 8'h07;
            16'd23942: data <= 8'hE0;
            16'd23943: data <= 8'h07;
            16'd23944: data <= 8'hE0;
            16'd23945: data <= 8'h07;
            16'd23946: data <= 8'hE0;
            16'd23947: data <= 8'h07;
            16'd23948: data <= 8'hE0;
            16'd23949: data <= 8'h07;
            16'd23950: data <= 8'hE0;
            16'd23951: data <= 8'h07;
            16'd23952: data <= 8'hE0;
            16'd23953: data <= 8'h07;
            16'd23954: data <= 8'hE0;
            16'd23955: data <= 8'h07;
            16'd23956: data <= 8'hE0;
            16'd23957: data <= 8'h07;
            16'd23958: data <= 8'hE0;
            16'd23959: data <= 8'h07;
            16'd23960: data <= 8'hFF;
            16'd23961: data <= 8'hFF;
            16'd23962: data <= 8'hE0;
            16'd23963: data <= 8'h07;
            16'd23964: data <= 8'hE0;
            16'd23965: data <= 8'h07;
            16'd23966: data <= 8'hE0;
            16'd23967: data <= 8'h07;
            16'd23968: data <= 8'hE0;
            16'd23969: data <= 8'h07;
            16'd23970: data <= 8'hE0;
            16'd23971: data <= 8'h07;
            16'd23972: data <= 8'hE0;
            16'd23973: data <= 8'h07;
            16'd23974: data <= 8'hE0;
            16'd23975: data <= 8'h07;
            16'd23976: data <= 8'hE0;
            16'd23977: data <= 8'h07;
            16'd23978: data <= 8'hE0;
            16'd23979: data <= 8'h07;
            16'd23980: data <= 8'hE0;
            16'd23981: data <= 8'h07;
            16'd23982: data <= 8'hE0;
            16'd23983: data <= 8'h07;
            16'd23984: data <= 8'hE0;
            16'd23985: data <= 8'h07;
            16'd23986: data <= 8'hE0;
            16'd23987: data <= 8'h07;
            16'd23988: data <= 8'hE0;
            16'd23989: data <= 8'h07;
            16'd23990: data <= 8'hE0;
            16'd23991: data <= 8'h07;
            16'd23992: data <= 8'hE0;
            16'd23993: data <= 8'h07;
            16'd23994: data <= 8'hE0;
            16'd23995: data <= 8'h07;
            16'd23996: data <= 8'hE0;
            16'd23997: data <= 8'h07;
            16'd23998: data <= 8'hE0;
            16'd23999: data <= 8'h07;
            16'd24000: data <= 8'hFF;
            16'd24001: data <= 8'hFF;
            16'd24002: data <= 8'hFF;
            16'd24003: data <= 8'hFF;
            16'd24004: data <= 8'hFF;
            16'd24005: data <= 8'hFF;
            16'd24006: data <= 8'hFF;
            16'd24007: data <= 8'hFF;
            16'd24008: data <= 8'hFF;
            16'd24009: data <= 8'hFF;
            16'd24010: data <= 8'hFF;
            16'd24011: data <= 8'hFF;
            16'd24012: data <= 8'hFF;
            16'd24013: data <= 8'hFF;
            16'd24014: data <= 8'hFF;
            16'd24015: data <= 8'hFF;
            16'd24016: data <= 8'hFF;
            16'd24017: data <= 8'hFF;
            16'd24018: data <= 8'hFF;
            16'd24019: data <= 8'hFF;
            16'd24020: data <= 8'hFF;
            16'd24021: data <= 8'hFF;
            16'd24022: data <= 8'hFF;
            16'd24023: data <= 8'hFF;
            16'd24024: data <= 8'hFF;
            16'd24025: data <= 8'hFF;
            16'd24026: data <= 8'hFF;
            16'd24027: data <= 8'hFF;
            16'd24028: data <= 8'hFF;
            16'd24029: data <= 8'hFF;
            16'd24030: data <= 8'hFF;
            16'd24031: data <= 8'hFF;
            16'd24032: data <= 8'hFF;
            16'd24033: data <= 8'hFF;
            16'd24034: data <= 8'hFF;
            16'd24035: data <= 8'hFF;
            16'd24036: data <= 8'hFF;
            16'd24037: data <= 8'hFF;
            16'd24038: data <= 8'hFF;
            16'd24039: data <= 8'hFF;
            16'd24040: data <= 8'hFF;
            16'd24041: data <= 8'hFF;
            16'd24042: data <= 8'hFF;
            16'd24043: data <= 8'hFF;
            16'd24044: data <= 8'hFF;
            16'd24045: data <= 8'hFF;
            16'd24046: data <= 8'hFF;
            16'd24047: data <= 8'hFF;
            16'd24048: data <= 8'hFF;
            16'd24049: data <= 8'hFF;
            16'd24050: data <= 8'hFF;
            16'd24051: data <= 8'hFF;
            16'd24052: data <= 8'hFF;
            16'd24053: data <= 8'hFF;
            16'd24054: data <= 8'hFF;
            16'd24055: data <= 8'hFF;
            16'd24056: data <= 8'hFF;
            16'd24057: data <= 8'hFF;
            16'd24058: data <= 8'hFF;
            16'd24059: data <= 8'hFF;
            16'd24060: data <= 8'hFF;
            16'd24061: data <= 8'hFF;
            16'd24062: data <= 8'hFF;
            16'd24063: data <= 8'hFF;
            16'd24064: data <= 8'hFF;
            16'd24065: data <= 8'hFF;
            16'd24066: data <= 8'hFF;
            16'd24067: data <= 8'hFF;
            16'd24068: data <= 8'hFF;
            16'd24069: data <= 8'hFF;
            16'd24070: data <= 8'hFF;
            16'd24071: data <= 8'hFF;
            16'd24072: data <= 8'hFF;
            16'd24073: data <= 8'hFF;
            16'd24074: data <= 8'hFF;
            16'd24075: data <= 8'hFF;
            16'd24076: data <= 8'hFF;
            16'd24077: data <= 8'hFF;
            16'd24078: data <= 8'hFF;
            16'd24079: data <= 8'hFF;
            16'd24080: data <= 8'hFF;
            16'd24081: data <= 8'hFF;
            16'd24082: data <= 8'hFF;
            16'd24083: data <= 8'hFF;
            16'd24084: data <= 8'hFF;
            16'd24085: data <= 8'hFF;
            16'd24086: data <= 8'hFF;
            16'd24087: data <= 8'hFF;
            16'd24088: data <= 8'hFF;
            16'd24089: data <= 8'hFF;
            16'd24090: data <= 8'hFF;
            16'd24091: data <= 8'hFF;
            16'd24092: data <= 8'hFF;
            16'd24093: data <= 8'hFF;
            16'd24094: data <= 8'hFF;
            16'd24095: data <= 8'hFF;
            16'd24096: data <= 8'hFF;
            16'd24097: data <= 8'hFF;
            16'd24098: data <= 8'hFF;
            16'd24099: data <= 8'hFF;
            16'd24100: data <= 8'hFF;
            16'd24101: data <= 8'hFF;
            16'd24102: data <= 8'hFF;
            16'd24103: data <= 8'hFF;
            16'd24104: data <= 8'hFF;
            16'd24105: data <= 8'hFF;
            16'd24106: data <= 8'hFF;
            16'd24107: data <= 8'hFF;
            16'd24108: data <= 8'hFF;
            16'd24109: data <= 8'hFF;
            16'd24110: data <= 8'hFF;
            16'd24111: data <= 8'hFF;
            16'd24112: data <= 8'hFF;
            16'd24113: data <= 8'hFF;
            16'd24114: data <= 8'hFF;
            16'd24115: data <= 8'hFF;
            16'd24116: data <= 8'hFF;
            16'd24117: data <= 8'hFF;
            16'd24118: data <= 8'hFF;
            16'd24119: data <= 8'hFF;
            16'd24120: data <= 8'hFF;
            16'd24121: data <= 8'hFF;
            16'd24122: data <= 8'hFF;
            16'd24123: data <= 8'hFF;
            16'd24124: data <= 8'hFF;
            16'd24125: data <= 8'hFF;
            16'd24126: data <= 8'hFF;
            16'd24127: data <= 8'hFF;
            16'd24128: data <= 8'hFF;
            16'd24129: data <= 8'hFF;
            16'd24130: data <= 8'hFF;
            16'd24131: data <= 8'hFF;
            16'd24132: data <= 8'hFF;
            16'd24133: data <= 8'hFF;
            16'd24134: data <= 8'hFF;
            16'd24135: data <= 8'hFF;
            16'd24136: data <= 8'hFF;
            16'd24137: data <= 8'hFF;
            16'd24138: data <= 8'hFF;
            16'd24139: data <= 8'hFF;
            16'd24140: data <= 8'hFF;
            16'd24141: data <= 8'hFF;
            16'd24142: data <= 8'hFF;
            16'd24143: data <= 8'hFF;
            16'd24144: data <= 8'hFF;
            16'd24145: data <= 8'hFF;
            16'd24146: data <= 8'hFF;
            16'd24147: data <= 8'hFF;
            16'd24148: data <= 8'hFF;
            16'd24149: data <= 8'hFF;
            16'd24150: data <= 8'hFF;
            16'd24151: data <= 8'hFF;
            16'd24152: data <= 8'hFF;
            16'd24153: data <= 8'hFF;
            16'd24154: data <= 8'hFF;
            16'd24155: data <= 8'hFF;
            16'd24156: data <= 8'hFF;
            16'd24157: data <= 8'hFF;
            16'd24158: data <= 8'hFF;
            16'd24159: data <= 8'hFF;
            16'd24160: data <= 8'hFF;
            16'd24161: data <= 8'hFF;
            16'd24162: data <= 8'hFF;
            16'd24163: data <= 8'hFF;
            16'd24164: data <= 8'hFF;
            16'd24165: data <= 8'hFF;
            16'd24166: data <= 8'hFF;
            16'd24167: data <= 8'hFF;
            16'd24168: data <= 8'hFF;
            16'd24169: data <= 8'hFF;
            16'd24170: data <= 8'hFF;
            16'd24171: data <= 8'hFF;
            16'd24172: data <= 8'hFF;
            16'd24173: data <= 8'hFF;
            16'd24174: data <= 8'hFF;
            16'd24175: data <= 8'hFF;
            16'd24176: data <= 8'hFF;
            16'd24177: data <= 8'hFF;
            16'd24178: data <= 8'hFF;
            16'd24179: data <= 8'hFF;
            16'd24180: data <= 8'hFF;
            16'd24181: data <= 8'hFF;
            16'd24182: data <= 8'hFF;
            16'd24183: data <= 8'hFF;
            16'd24184: data <= 8'hFF;
            16'd24185: data <= 8'hFF;
            16'd24186: data <= 8'hFF;
            16'd24187: data <= 8'hFF;
            16'd24188: data <= 8'hFF;
            16'd24189: data <= 8'hFF;
            16'd24190: data <= 8'hFF;
            16'd24191: data <= 8'hFF;
            16'd24192: data <= 8'hFF;
            16'd24193: data <= 8'hFF;
            16'd24194: data <= 8'hFF;
            16'd24195: data <= 8'hFF;
            16'd24196: data <= 8'hFF;
            16'd24197: data <= 8'hFF;
            16'd24198: data <= 8'hFF;
            16'd24199: data <= 8'hFF;
            16'd24200: data <= 8'hFF;
            16'd24201: data <= 8'hFF;
            16'd24202: data <= 8'hFF;
            16'd24203: data <= 8'hFF;
            16'd24204: data <= 8'hFF;
            16'd24205: data <= 8'hFF;
            16'd24206: data <= 8'hFF;
            16'd24207: data <= 8'hFF;
            16'd24208: data <= 8'hFF;
            16'd24209: data <= 8'hFF;
            16'd24210: data <= 8'hFF;
            16'd24211: data <= 8'hFF;
            16'd24212: data <= 8'hFF;
            16'd24213: data <= 8'hFF;
            16'd24214: data <= 8'hFF;
            16'd24215: data <= 8'hFF;
            16'd24216: data <= 8'hFF;
            16'd24217: data <= 8'hFF;
            16'd24218: data <= 8'hFF;
            16'd24219: data <= 8'hFF;
            16'd24220: data <= 8'hFF;
            16'd24221: data <= 8'hFF;
            16'd24222: data <= 8'hFF;
            16'd24223: data <= 8'hFF;
            16'd24224: data <= 8'hFF;
            16'd24225: data <= 8'hFF;
            16'd24226: data <= 8'hFF;
            16'd24227: data <= 8'hFF;
            16'd24228: data <= 8'hFF;
            16'd24229: data <= 8'hFF;
            16'd24230: data <= 8'hFF;
            16'd24231: data <= 8'hFF;
            16'd24232: data <= 8'hFF;
            16'd24233: data <= 8'hFF;
            16'd24234: data <= 8'hFF;
            16'd24235: data <= 8'hFF;
            16'd24236: data <= 8'hFF;
            16'd24237: data <= 8'hFF;
            16'd24238: data <= 8'hFF;
            16'd24239: data <= 8'hFF;
            16'd24240: data <= 8'hFF;
            16'd24241: data <= 8'hFF;
            16'd24242: data <= 8'hE0;
            16'd24243: data <= 8'h07;
            16'd24244: data <= 8'hE0;
            16'd24245: data <= 8'h07;
            16'd24246: data <= 8'hE0;
            16'd24247: data <= 8'h07;
            16'd24248: data <= 8'hE0;
            16'd24249: data <= 8'h07;
            16'd24250: data <= 8'hE0;
            16'd24251: data <= 8'h07;
            16'd24252: data <= 8'hE0;
            16'd24253: data <= 8'h07;
            16'd24254: data <= 8'hE0;
            16'd24255: data <= 8'h07;
            16'd24256: data <= 8'hE0;
            16'd24257: data <= 8'h07;
            16'd24258: data <= 8'hE0;
            16'd24259: data <= 8'h07;
            16'd24260: data <= 8'hE0;
            16'd24261: data <= 8'h07;
            16'd24262: data <= 8'hE0;
            16'd24263: data <= 8'h07;
            16'd24264: data <= 8'hE0;
            16'd24265: data <= 8'h07;
            16'd24266: data <= 8'hE0;
            16'd24267: data <= 8'h07;
            16'd24268: data <= 8'hE0;
            16'd24269: data <= 8'h07;
            16'd24270: data <= 8'hE0;
            16'd24271: data <= 8'h07;
            16'd24272: data <= 8'hE0;
            16'd24273: data <= 8'h07;
            16'd24274: data <= 8'hE0;
            16'd24275: data <= 8'h07;
            16'd24276: data <= 8'hE0;
            16'd24277: data <= 8'h07;
            16'd24278: data <= 8'hE0;
            16'd24279: data <= 8'h07;
            16'd24280: data <= 8'hFF;
            16'd24281: data <= 8'hFF;
            16'd24282: data <= 8'hE0;
            16'd24283: data <= 8'h07;
            16'd24284: data <= 8'hE0;
            16'd24285: data <= 8'h07;
            16'd24286: data <= 8'hE0;
            16'd24287: data <= 8'h07;
            16'd24288: data <= 8'hE0;
            16'd24289: data <= 8'h07;
            16'd24290: data <= 8'hE0;
            16'd24291: data <= 8'h07;
            16'd24292: data <= 8'hE0;
            16'd24293: data <= 8'h07;
            16'd24294: data <= 8'hE0;
            16'd24295: data <= 8'h07;
            16'd24296: data <= 8'hE0;
            16'd24297: data <= 8'h07;
            16'd24298: data <= 8'hE0;
            16'd24299: data <= 8'h07;
            16'd24300: data <= 8'hE0;
            16'd24301: data <= 8'h07;
            16'd24302: data <= 8'hE0;
            16'd24303: data <= 8'h07;
            16'd24304: data <= 8'hE0;
            16'd24305: data <= 8'h07;
            16'd24306: data <= 8'hE0;
            16'd24307: data <= 8'h07;
            16'd24308: data <= 8'hE0;
            16'd24309: data <= 8'h07;
            16'd24310: data <= 8'hE0;
            16'd24311: data <= 8'h07;
            16'd24312: data <= 8'hE0;
            16'd24313: data <= 8'h07;
            16'd24314: data <= 8'hE0;
            16'd24315: data <= 8'h07;
            16'd24316: data <= 8'hE0;
            16'd24317: data <= 8'h07;
            16'd24318: data <= 8'hE0;
            16'd24319: data <= 8'h07;
            16'd24320: data <= 8'hFF;
            16'd24321: data <= 8'hFF;
            16'd24322: data <= 8'hE0;
            16'd24323: data <= 8'h07;
            16'd24324: data <= 8'hE0;
            16'd24325: data <= 8'h07;
            16'd24326: data <= 8'hE0;
            16'd24327: data <= 8'h07;
            16'd24328: data <= 8'hE0;
            16'd24329: data <= 8'h07;
            16'd24330: data <= 8'hE0;
            16'd24331: data <= 8'h07;
            16'd24332: data <= 8'hE0;
            16'd24333: data <= 8'h07;
            16'd24334: data <= 8'hE0;
            16'd24335: data <= 8'h07;
            16'd24336: data <= 8'hE0;
            16'd24337: data <= 8'h07;
            16'd24338: data <= 8'hE0;
            16'd24339: data <= 8'h07;
            16'd24340: data <= 8'hE0;
            16'd24341: data <= 8'h07;
            16'd24342: data <= 8'hE0;
            16'd24343: data <= 8'h07;
            16'd24344: data <= 8'hE0;
            16'd24345: data <= 8'h07;
            16'd24346: data <= 8'hE0;
            16'd24347: data <= 8'h07;
            16'd24348: data <= 8'hE0;
            16'd24349: data <= 8'h07;
            16'd24350: data <= 8'hE0;
            16'd24351: data <= 8'h07;
            16'd24352: data <= 8'hE0;
            16'd24353: data <= 8'h07;
            16'd24354: data <= 8'hE0;
            16'd24355: data <= 8'h07;
            16'd24356: data <= 8'hE0;
            16'd24357: data <= 8'h07;
            16'd24358: data <= 8'hE0;
            16'd24359: data <= 8'h07;
            16'd24360: data <= 8'hFF;
            16'd24361: data <= 8'hFF;
            16'd24362: data <= 8'hE0;
            16'd24363: data <= 8'h07;
            16'd24364: data <= 8'hE0;
            16'd24365: data <= 8'h07;
            16'd24366: data <= 8'hE0;
            16'd24367: data <= 8'h07;
            16'd24368: data <= 8'hE0;
            16'd24369: data <= 8'h07;
            16'd24370: data <= 8'hE0;
            16'd24371: data <= 8'h07;
            16'd24372: data <= 8'hE0;
            16'd24373: data <= 8'h07;
            16'd24374: data <= 8'hE0;
            16'd24375: data <= 8'h07;
            16'd24376: data <= 8'hE0;
            16'd24377: data <= 8'h07;
            16'd24378: data <= 8'hE0;
            16'd24379: data <= 8'h07;
            16'd24380: data <= 8'hE0;
            16'd24381: data <= 8'h07;
            16'd24382: data <= 8'hE0;
            16'd24383: data <= 8'h07;
            16'd24384: data <= 8'hE0;
            16'd24385: data <= 8'h07;
            16'd24386: data <= 8'hE0;
            16'd24387: data <= 8'h07;
            16'd24388: data <= 8'hE0;
            16'd24389: data <= 8'h07;
            16'd24390: data <= 8'hE0;
            16'd24391: data <= 8'h07;
            16'd24392: data <= 8'hE0;
            16'd24393: data <= 8'h07;
            16'd24394: data <= 8'hE0;
            16'd24395: data <= 8'h07;
            16'd24396: data <= 8'hE0;
            16'd24397: data <= 8'h07;
            16'd24398: data <= 8'hE0;
            16'd24399: data <= 8'h07;
            16'd24400: data <= 8'hFF;
            16'd24401: data <= 8'hFF;
            16'd24402: data <= 8'hE0;
            16'd24403: data <= 8'h07;
            16'd24404: data <= 8'hE0;
            16'd24405: data <= 8'h07;
            16'd24406: data <= 8'hE0;
            16'd24407: data <= 8'h07;
            16'd24408: data <= 8'hE0;
            16'd24409: data <= 8'h07;
            16'd24410: data <= 8'hE0;
            16'd24411: data <= 8'h07;
            16'd24412: data <= 8'hE0;
            16'd24413: data <= 8'h07;
            16'd24414: data <= 8'hE0;
            16'd24415: data <= 8'h07;
            16'd24416: data <= 8'hE0;
            16'd24417: data <= 8'h07;
            16'd24418: data <= 8'hE0;
            16'd24419: data <= 8'h07;
            16'd24420: data <= 8'hE0;
            16'd24421: data <= 8'h07;
            16'd24422: data <= 8'hE0;
            16'd24423: data <= 8'h07;
            16'd24424: data <= 8'hE0;
            16'd24425: data <= 8'h07;
            16'd24426: data <= 8'hE0;
            16'd24427: data <= 8'h07;
            16'd24428: data <= 8'hE0;
            16'd24429: data <= 8'h07;
            16'd24430: data <= 8'hE0;
            16'd24431: data <= 8'h07;
            16'd24432: data <= 8'hE0;
            16'd24433: data <= 8'h07;
            16'd24434: data <= 8'hE0;
            16'd24435: data <= 8'h07;
            16'd24436: data <= 8'hE0;
            16'd24437: data <= 8'h07;
            16'd24438: data <= 8'hE0;
            16'd24439: data <= 8'h07;
            16'd24440: data <= 8'hFF;
            16'd24441: data <= 8'hFF;
            16'd24442: data <= 8'hE0;
            16'd24443: data <= 8'h07;
            16'd24444: data <= 8'hE0;
            16'd24445: data <= 8'h07;
            16'd24446: data <= 8'hE0;
            16'd24447: data <= 8'h07;
            16'd24448: data <= 8'hE0;
            16'd24449: data <= 8'h07;
            16'd24450: data <= 8'hE0;
            16'd24451: data <= 8'h07;
            16'd24452: data <= 8'hE0;
            16'd24453: data <= 8'h07;
            16'd24454: data <= 8'hE0;
            16'd24455: data <= 8'h07;
            16'd24456: data <= 8'hE0;
            16'd24457: data <= 8'h07;
            16'd24458: data <= 8'hE0;
            16'd24459: data <= 8'h07;
            16'd24460: data <= 8'hE0;
            16'd24461: data <= 8'h07;
            16'd24462: data <= 8'hE0;
            16'd24463: data <= 8'h07;
            16'd24464: data <= 8'hE0;
            16'd24465: data <= 8'h07;
            16'd24466: data <= 8'hE0;
            16'd24467: data <= 8'h07;
            16'd24468: data <= 8'hE0;
            16'd24469: data <= 8'h07;
            16'd24470: data <= 8'hE0;
            16'd24471: data <= 8'h07;
            16'd24472: data <= 8'hE0;
            16'd24473: data <= 8'h07;
            16'd24474: data <= 8'hE0;
            16'd24475: data <= 8'h07;
            16'd24476: data <= 8'hE0;
            16'd24477: data <= 8'h07;
            16'd24478: data <= 8'hE0;
            16'd24479: data <= 8'h07;
            16'd24480: data <= 8'hFF;
            16'd24481: data <= 8'hFF;
            16'd24482: data <= 8'hE0;
            16'd24483: data <= 8'h07;
            16'd24484: data <= 8'hE0;
            16'd24485: data <= 8'h07;
            16'd24486: data <= 8'hE0;
            16'd24487: data <= 8'h07;
            16'd24488: data <= 8'hE0;
            16'd24489: data <= 8'h07;
            16'd24490: data <= 8'hE0;
            16'd24491: data <= 8'h07;
            16'd24492: data <= 8'hE0;
            16'd24493: data <= 8'h07;
            16'd24494: data <= 8'hE0;
            16'd24495: data <= 8'h07;
            16'd24496: data <= 8'hE0;
            16'd24497: data <= 8'h07;
            16'd24498: data <= 8'hE0;
            16'd24499: data <= 8'h07;
            16'd24500: data <= 8'hE0;
            16'd24501: data <= 8'h07;
            16'd24502: data <= 8'hE0;
            16'd24503: data <= 8'h07;
            16'd24504: data <= 8'hE0;
            16'd24505: data <= 8'h07;
            16'd24506: data <= 8'hE0;
            16'd24507: data <= 8'h07;
            16'd24508: data <= 8'hE0;
            16'd24509: data <= 8'h07;
            16'd24510: data <= 8'hE0;
            16'd24511: data <= 8'h07;
            16'd24512: data <= 8'hE0;
            16'd24513: data <= 8'h07;
            16'd24514: data <= 8'hE0;
            16'd24515: data <= 8'h07;
            16'd24516: data <= 8'hE0;
            16'd24517: data <= 8'h07;
            16'd24518: data <= 8'hE0;
            16'd24519: data <= 8'h07;
            16'd24520: data <= 8'hFF;
            16'd24521: data <= 8'hFF;
            16'd24522: data <= 8'hE0;
            16'd24523: data <= 8'h07;
            16'd24524: data <= 8'hE0;
            16'd24525: data <= 8'h07;
            16'd24526: data <= 8'hE0;
            16'd24527: data <= 8'h07;
            16'd24528: data <= 8'hE0;
            16'd24529: data <= 8'h07;
            16'd24530: data <= 8'hE0;
            16'd24531: data <= 8'h07;
            16'd24532: data <= 8'hE0;
            16'd24533: data <= 8'h07;
            16'd24534: data <= 8'hE0;
            16'd24535: data <= 8'h07;
            16'd24536: data <= 8'hE0;
            16'd24537: data <= 8'h07;
            16'd24538: data <= 8'hE0;
            16'd24539: data <= 8'h07;
            16'd24540: data <= 8'hE0;
            16'd24541: data <= 8'h07;
            16'd24542: data <= 8'hE0;
            16'd24543: data <= 8'h07;
            16'd24544: data <= 8'hE0;
            16'd24545: data <= 8'h07;
            16'd24546: data <= 8'hE0;
            16'd24547: data <= 8'h07;
            16'd24548: data <= 8'hE0;
            16'd24549: data <= 8'h07;
            16'd24550: data <= 8'hE0;
            16'd24551: data <= 8'h07;
            16'd24552: data <= 8'hE0;
            16'd24553: data <= 8'h07;
            16'd24554: data <= 8'hE0;
            16'd24555: data <= 8'h07;
            16'd24556: data <= 8'hE0;
            16'd24557: data <= 8'h07;
            16'd24558: data <= 8'hE0;
            16'd24559: data <= 8'h07;
            16'd24560: data <= 8'hFF;
            16'd24561: data <= 8'hFF;
            16'd24562: data <= 8'hE0;
            16'd24563: data <= 8'h07;
            16'd24564: data <= 8'hE0;
            16'd24565: data <= 8'h07;
            16'd24566: data <= 8'hE0;
            16'd24567: data <= 8'h07;
            16'd24568: data <= 8'hE0;
            16'd24569: data <= 8'h07;
            16'd24570: data <= 8'hE0;
            16'd24571: data <= 8'h07;
            16'd24572: data <= 8'hE0;
            16'd24573: data <= 8'h07;
            16'd24574: data <= 8'hE0;
            16'd24575: data <= 8'h07;
            16'd24576: data <= 8'hE0;
            16'd24577: data <= 8'h07;
            16'd24578: data <= 8'hE0;
            16'd24579: data <= 8'h07;
            16'd24580: data <= 8'hE0;
            16'd24581: data <= 8'h07;
            16'd24582: data <= 8'hE0;
            16'd24583: data <= 8'h07;
            16'd24584: data <= 8'hE0;
            16'd24585: data <= 8'h07;
            16'd24586: data <= 8'hE0;
            16'd24587: data <= 8'h07;
            16'd24588: data <= 8'hE0;
            16'd24589: data <= 8'h07;
            16'd24590: data <= 8'hE0;
            16'd24591: data <= 8'h07;
            16'd24592: data <= 8'hE0;
            16'd24593: data <= 8'h07;
            16'd24594: data <= 8'hE0;
            16'd24595: data <= 8'h07;
            16'd24596: data <= 8'hE0;
            16'd24597: data <= 8'h07;
            16'd24598: data <= 8'hE0;
            16'd24599: data <= 8'h07;
            16'd24600: data <= 8'hFF;
            16'd24601: data <= 8'hFF;
            16'd24602: data <= 8'hE0;
            16'd24603: data <= 8'h07;
            16'd24604: data <= 8'hE0;
            16'd24605: data <= 8'h07;
            16'd24606: data <= 8'hE0;
            16'd24607: data <= 8'h07;
            16'd24608: data <= 8'hE0;
            16'd24609: data <= 8'h07;
            16'd24610: data <= 8'hE0;
            16'd24611: data <= 8'h07;
            16'd24612: data <= 8'hE0;
            16'd24613: data <= 8'h07;
            16'd24614: data <= 8'hE0;
            16'd24615: data <= 8'h07;
            16'd24616: data <= 8'hE0;
            16'd24617: data <= 8'h07;
            16'd24618: data <= 8'hE0;
            16'd24619: data <= 8'h07;
            16'd24620: data <= 8'hE0;
            16'd24621: data <= 8'h07;
            16'd24622: data <= 8'hE0;
            16'd24623: data <= 8'h07;
            16'd24624: data <= 8'hE0;
            16'd24625: data <= 8'h07;
            16'd24626: data <= 8'hE0;
            16'd24627: data <= 8'h07;
            16'd24628: data <= 8'hE0;
            16'd24629: data <= 8'h07;
            16'd24630: data <= 8'hE0;
            16'd24631: data <= 8'h07;
            16'd24632: data <= 8'hE0;
            16'd24633: data <= 8'h07;
            16'd24634: data <= 8'hE0;
            16'd24635: data <= 8'h07;
            16'd24636: data <= 8'hE0;
            16'd24637: data <= 8'h07;
            16'd24638: data <= 8'hE0;
            16'd24639: data <= 8'h07;
            16'd24640: data <= 8'hFF;
            16'd24641: data <= 8'hFF;
            16'd24642: data <= 8'hE0;
            16'd24643: data <= 8'h07;
            16'd24644: data <= 8'hE0;
            16'd24645: data <= 8'h07;
            16'd24646: data <= 8'hE0;
            16'd24647: data <= 8'h07;
            16'd24648: data <= 8'hE0;
            16'd24649: data <= 8'h07;
            16'd24650: data <= 8'hE0;
            16'd24651: data <= 8'h07;
            16'd24652: data <= 8'hE0;
            16'd24653: data <= 8'h07;
            16'd24654: data <= 8'hE0;
            16'd24655: data <= 8'h07;
            16'd24656: data <= 8'hE0;
            16'd24657: data <= 8'h07;
            16'd24658: data <= 8'hE0;
            16'd24659: data <= 8'h07;
            16'd24660: data <= 8'hE0;
            16'd24661: data <= 8'h07;
            16'd24662: data <= 8'hE0;
            16'd24663: data <= 8'h07;
            16'd24664: data <= 8'hE0;
            16'd24665: data <= 8'h07;
            16'd24666: data <= 8'hE0;
            16'd24667: data <= 8'h07;
            16'd24668: data <= 8'hE0;
            16'd24669: data <= 8'h07;
            16'd24670: data <= 8'hE0;
            16'd24671: data <= 8'h07;
            16'd24672: data <= 8'hE0;
            16'd24673: data <= 8'h07;
            16'd24674: data <= 8'hE0;
            16'd24675: data <= 8'h07;
            16'd24676: data <= 8'hE0;
            16'd24677: data <= 8'h07;
            16'd24678: data <= 8'hE0;
            16'd24679: data <= 8'h07;
            16'd24680: data <= 8'hFF;
            16'd24681: data <= 8'hFF;
            16'd24682: data <= 8'hE0;
            16'd24683: data <= 8'h07;
            16'd24684: data <= 8'hE0;
            16'd24685: data <= 8'h07;
            16'd24686: data <= 8'hE0;
            16'd24687: data <= 8'h07;
            16'd24688: data <= 8'hE0;
            16'd24689: data <= 8'h07;
            16'd24690: data <= 8'hE0;
            16'd24691: data <= 8'h07;
            16'd24692: data <= 8'hE0;
            16'd24693: data <= 8'h07;
            16'd24694: data <= 8'hE0;
            16'd24695: data <= 8'h07;
            16'd24696: data <= 8'hE0;
            16'd24697: data <= 8'h07;
            16'd24698: data <= 8'hE0;
            16'd24699: data <= 8'h07;
            16'd24700: data <= 8'hE0;
            16'd24701: data <= 8'h07;
            16'd24702: data <= 8'hE0;
            16'd24703: data <= 8'h07;
            16'd24704: data <= 8'hE0;
            16'd24705: data <= 8'h07;
            16'd24706: data <= 8'hE0;
            16'd24707: data <= 8'h07;
            16'd24708: data <= 8'hE0;
            16'd24709: data <= 8'h07;
            16'd24710: data <= 8'hE0;
            16'd24711: data <= 8'h07;
            16'd24712: data <= 8'hE0;
            16'd24713: data <= 8'h07;
            16'd24714: data <= 8'hE0;
            16'd24715: data <= 8'h07;
            16'd24716: data <= 8'hE0;
            16'd24717: data <= 8'h07;
            16'd24718: data <= 8'hE0;
            16'd24719: data <= 8'h07;
            16'd24720: data <= 8'hFF;
            16'd24721: data <= 8'hFF;
            16'd24722: data <= 8'hE0;
            16'd24723: data <= 8'h07;
            16'd24724: data <= 8'hE0;
            16'd24725: data <= 8'h07;
            16'd24726: data <= 8'hE0;
            16'd24727: data <= 8'h07;
            16'd24728: data <= 8'hE0;
            16'd24729: data <= 8'h07;
            16'd24730: data <= 8'hE0;
            16'd24731: data <= 8'h07;
            16'd24732: data <= 8'hE0;
            16'd24733: data <= 8'h07;
            16'd24734: data <= 8'hE0;
            16'd24735: data <= 8'h07;
            16'd24736: data <= 8'hE0;
            16'd24737: data <= 8'h07;
            16'd24738: data <= 8'hE0;
            16'd24739: data <= 8'h07;
            16'd24740: data <= 8'hE0;
            16'd24741: data <= 8'h07;
            16'd24742: data <= 8'hE0;
            16'd24743: data <= 8'h07;
            16'd24744: data <= 8'hE0;
            16'd24745: data <= 8'h07;
            16'd24746: data <= 8'hE0;
            16'd24747: data <= 8'h07;
            16'd24748: data <= 8'hE0;
            16'd24749: data <= 8'h07;
            16'd24750: data <= 8'hE0;
            16'd24751: data <= 8'h07;
            16'd24752: data <= 8'hE0;
            16'd24753: data <= 8'h07;
            16'd24754: data <= 8'hE0;
            16'd24755: data <= 8'h07;
            16'd24756: data <= 8'hE0;
            16'd24757: data <= 8'h07;
            16'd24758: data <= 8'hE0;
            16'd24759: data <= 8'h07;
            16'd24760: data <= 8'hFF;
            16'd24761: data <= 8'hFF;
            16'd24762: data <= 8'hE0;
            16'd24763: data <= 8'h07;
            16'd24764: data <= 8'hE0;
            16'd24765: data <= 8'h07;
            16'd24766: data <= 8'hE0;
            16'd24767: data <= 8'h07;
            16'd24768: data <= 8'hE0;
            16'd24769: data <= 8'h07;
            16'd24770: data <= 8'hE0;
            16'd24771: data <= 8'h07;
            16'd24772: data <= 8'hE0;
            16'd24773: data <= 8'h07;
            16'd24774: data <= 8'hE0;
            16'd24775: data <= 8'h07;
            16'd24776: data <= 8'hE0;
            16'd24777: data <= 8'h07;
            16'd24778: data <= 8'hE0;
            16'd24779: data <= 8'h07;
            16'd24780: data <= 8'hE0;
            16'd24781: data <= 8'h07;
            16'd24782: data <= 8'hE0;
            16'd24783: data <= 8'h07;
            16'd24784: data <= 8'hE0;
            16'd24785: data <= 8'h07;
            16'd24786: data <= 8'hE0;
            16'd24787: data <= 8'h07;
            16'd24788: data <= 8'hE0;
            16'd24789: data <= 8'h07;
            16'd24790: data <= 8'hE0;
            16'd24791: data <= 8'h07;
            16'd24792: data <= 8'hE0;
            16'd24793: data <= 8'h07;
            16'd24794: data <= 8'hE0;
            16'd24795: data <= 8'h07;
            16'd24796: data <= 8'hE0;
            16'd24797: data <= 8'h07;
            16'd24798: data <= 8'hE0;
            16'd24799: data <= 8'h07;
            16'd24800: data <= 8'hFF;
            16'd24801: data <= 8'hFF;
            16'd24802: data <= 8'hE0;
            16'd24803: data <= 8'h07;
            16'd24804: data <= 8'hE0;
            16'd24805: data <= 8'h07;
            16'd24806: data <= 8'hE0;
            16'd24807: data <= 8'h07;
            16'd24808: data <= 8'hE0;
            16'd24809: data <= 8'h07;
            16'd24810: data <= 8'hE0;
            16'd24811: data <= 8'h07;
            16'd24812: data <= 8'hE0;
            16'd24813: data <= 8'h07;
            16'd24814: data <= 8'hE0;
            16'd24815: data <= 8'h07;
            16'd24816: data <= 8'hE0;
            16'd24817: data <= 8'h07;
            16'd24818: data <= 8'hE0;
            16'd24819: data <= 8'h07;
            16'd24820: data <= 8'hE0;
            16'd24821: data <= 8'h07;
            16'd24822: data <= 8'hE0;
            16'd24823: data <= 8'h07;
            16'd24824: data <= 8'hE0;
            16'd24825: data <= 8'h07;
            16'd24826: data <= 8'hE0;
            16'd24827: data <= 8'h07;
            16'd24828: data <= 8'hE0;
            16'd24829: data <= 8'h07;
            16'd24830: data <= 8'hE0;
            16'd24831: data <= 8'h07;
            16'd24832: data <= 8'hE0;
            16'd24833: data <= 8'h07;
            16'd24834: data <= 8'hE0;
            16'd24835: data <= 8'h07;
            16'd24836: data <= 8'hE0;
            16'd24837: data <= 8'h07;
            16'd24838: data <= 8'hE0;
            16'd24839: data <= 8'h07;
            16'd24840: data <= 8'hFF;
            16'd24841: data <= 8'hFF;
            16'd24842: data <= 8'hE0;
            16'd24843: data <= 8'h07;
            16'd24844: data <= 8'hE0;
            16'd24845: data <= 8'h07;
            16'd24846: data <= 8'hE0;
            16'd24847: data <= 8'h07;
            16'd24848: data <= 8'hE0;
            16'd24849: data <= 8'h07;
            16'd24850: data <= 8'hE0;
            16'd24851: data <= 8'h07;
            16'd24852: data <= 8'hE0;
            16'd24853: data <= 8'h07;
            16'd24854: data <= 8'hE0;
            16'd24855: data <= 8'h07;
            16'd24856: data <= 8'hE0;
            16'd24857: data <= 8'h07;
            16'd24858: data <= 8'hE0;
            16'd24859: data <= 8'h07;
            16'd24860: data <= 8'hE0;
            16'd24861: data <= 8'h07;
            16'd24862: data <= 8'hE0;
            16'd24863: data <= 8'h07;
            16'd24864: data <= 8'hE0;
            16'd24865: data <= 8'h07;
            16'd24866: data <= 8'hE0;
            16'd24867: data <= 8'h07;
            16'd24868: data <= 8'hE0;
            16'd24869: data <= 8'h07;
            16'd24870: data <= 8'hE0;
            16'd24871: data <= 8'h07;
            16'd24872: data <= 8'hE0;
            16'd24873: data <= 8'h07;
            16'd24874: data <= 8'hE0;
            16'd24875: data <= 8'h07;
            16'd24876: data <= 8'hE0;
            16'd24877: data <= 8'h07;
            16'd24878: data <= 8'hE0;
            16'd24879: data <= 8'h07;
            16'd24880: data <= 8'hFF;
            16'd24881: data <= 8'hFF;
            16'd24882: data <= 8'hE0;
            16'd24883: data <= 8'h07;
            16'd24884: data <= 8'hE0;
            16'd24885: data <= 8'h07;
            16'd24886: data <= 8'hE0;
            16'd24887: data <= 8'h07;
            16'd24888: data <= 8'hE0;
            16'd24889: data <= 8'h07;
            16'd24890: data <= 8'hE0;
            16'd24891: data <= 8'h07;
            16'd24892: data <= 8'hE0;
            16'd24893: data <= 8'h07;
            16'd24894: data <= 8'hE0;
            16'd24895: data <= 8'h07;
            16'd24896: data <= 8'hE0;
            16'd24897: data <= 8'h07;
            16'd24898: data <= 8'hE0;
            16'd24899: data <= 8'h07;
            16'd24900: data <= 8'hE0;
            16'd24901: data <= 8'h07;
            16'd24902: data <= 8'hE0;
            16'd24903: data <= 8'h07;
            16'd24904: data <= 8'hE0;
            16'd24905: data <= 8'h07;
            16'd24906: data <= 8'hE0;
            16'd24907: data <= 8'h07;
            16'd24908: data <= 8'hE0;
            16'd24909: data <= 8'h07;
            16'd24910: data <= 8'hE0;
            16'd24911: data <= 8'h07;
            16'd24912: data <= 8'hE0;
            16'd24913: data <= 8'h07;
            16'd24914: data <= 8'hE0;
            16'd24915: data <= 8'h07;
            16'd24916: data <= 8'hE0;
            16'd24917: data <= 8'h07;
            16'd24918: data <= 8'hE0;
            16'd24919: data <= 8'h07;
            16'd24920: data <= 8'hFF;
            16'd24921: data <= 8'hFF;
            16'd24922: data <= 8'hE0;
            16'd24923: data <= 8'h07;
            16'd24924: data <= 8'hE0;
            16'd24925: data <= 8'h07;
            16'd24926: data <= 8'hE0;
            16'd24927: data <= 8'h07;
            16'd24928: data <= 8'hE0;
            16'd24929: data <= 8'h07;
            16'd24930: data <= 8'hE0;
            16'd24931: data <= 8'h07;
            16'd24932: data <= 8'hE0;
            16'd24933: data <= 8'h07;
            16'd24934: data <= 8'hE0;
            16'd24935: data <= 8'h07;
            16'd24936: data <= 8'hE0;
            16'd24937: data <= 8'h07;
            16'd24938: data <= 8'hE0;
            16'd24939: data <= 8'h07;
            16'd24940: data <= 8'hE0;
            16'd24941: data <= 8'h07;
            16'd24942: data <= 8'hE0;
            16'd24943: data <= 8'h07;
            16'd24944: data <= 8'hE0;
            16'd24945: data <= 8'h07;
            16'd24946: data <= 8'hE0;
            16'd24947: data <= 8'h07;
            16'd24948: data <= 8'hE0;
            16'd24949: data <= 8'h07;
            16'd24950: data <= 8'hE0;
            16'd24951: data <= 8'h07;
            16'd24952: data <= 8'hE0;
            16'd24953: data <= 8'h07;
            16'd24954: data <= 8'hE0;
            16'd24955: data <= 8'h07;
            16'd24956: data <= 8'hE0;
            16'd24957: data <= 8'h07;
            16'd24958: data <= 8'hE0;
            16'd24959: data <= 8'h07;
            16'd24960: data <= 8'hFF;
            16'd24961: data <= 8'hFF;
            16'd24962: data <= 8'hE0;
            16'd24963: data <= 8'h07;
            16'd24964: data <= 8'hE0;
            16'd24965: data <= 8'h07;
            16'd24966: data <= 8'hE0;
            16'd24967: data <= 8'h07;
            16'd24968: data <= 8'hE0;
            16'd24969: data <= 8'h07;
            16'd24970: data <= 8'hE0;
            16'd24971: data <= 8'h07;
            16'd24972: data <= 8'hE0;
            16'd24973: data <= 8'h07;
            16'd24974: data <= 8'hE0;
            16'd24975: data <= 8'h07;
            16'd24976: data <= 8'hE0;
            16'd24977: data <= 8'h07;
            16'd24978: data <= 8'hE0;
            16'd24979: data <= 8'h07;
            16'd24980: data <= 8'hE0;
            16'd24981: data <= 8'h07;
            16'd24982: data <= 8'hE0;
            16'd24983: data <= 8'h07;
            16'd24984: data <= 8'hE0;
            16'd24985: data <= 8'h07;
            16'd24986: data <= 8'hE0;
            16'd24987: data <= 8'h07;
            16'd24988: data <= 8'hE0;
            16'd24989: data <= 8'h07;
            16'd24990: data <= 8'hE0;
            16'd24991: data <= 8'h07;
            16'd24992: data <= 8'hE0;
            16'd24993: data <= 8'h07;
            16'd24994: data <= 8'hE0;
            16'd24995: data <= 8'h07;
            16'd24996: data <= 8'hE0;
            16'd24997: data <= 8'h07;
            16'd24998: data <= 8'hE0;
            16'd24999: data <= 8'h07;
            16'd25000: data <= 8'hFF;
            16'd25001: data <= 8'hFF;
            16'd25002: data <= 8'hE0;
            16'd25003: data <= 8'h07;
            16'd25004: data <= 8'hE0;
            16'd25005: data <= 8'h07;
            16'd25006: data <= 8'hE0;
            16'd25007: data <= 8'h07;
            16'd25008: data <= 8'hE0;
            16'd25009: data <= 8'h07;
            16'd25010: data <= 8'hE0;
            16'd25011: data <= 8'h07;
            16'd25012: data <= 8'hE0;
            16'd25013: data <= 8'h07;
            16'd25014: data <= 8'hE0;
            16'd25015: data <= 8'h07;
            16'd25016: data <= 8'hE0;
            16'd25017: data <= 8'h07;
            16'd25018: data <= 8'hE0;
            16'd25019: data <= 8'h07;
            16'd25020: data <= 8'hE0;
            16'd25021: data <= 8'h07;
            16'd25022: data <= 8'hE0;
            16'd25023: data <= 8'h07;
            16'd25024: data <= 8'hE0;
            16'd25025: data <= 8'h07;
            16'd25026: data <= 8'hE0;
            16'd25027: data <= 8'h07;
            16'd25028: data <= 8'hE0;
            16'd25029: data <= 8'h07;
            16'd25030: data <= 8'hE0;
            16'd25031: data <= 8'h07;
            16'd25032: data <= 8'hE0;
            16'd25033: data <= 8'h07;
            16'd25034: data <= 8'hE0;
            16'd25035: data <= 8'h07;
            16'd25036: data <= 8'hE0;
            16'd25037: data <= 8'h07;
            16'd25038: data <= 8'hE0;
            16'd25039: data <= 8'h07;
            16'd25040: data <= 8'hFF;
            16'd25041: data <= 8'hFF;
            16'd25042: data <= 8'hE0;
            16'd25043: data <= 8'h07;
            16'd25044: data <= 8'hE0;
            16'd25045: data <= 8'h07;
            16'd25046: data <= 8'hE0;
            16'd25047: data <= 8'h07;
            16'd25048: data <= 8'hE0;
            16'd25049: data <= 8'h07;
            16'd25050: data <= 8'hE0;
            16'd25051: data <= 8'h07;
            16'd25052: data <= 8'hE0;
            16'd25053: data <= 8'h07;
            16'd25054: data <= 8'hE0;
            16'd25055: data <= 8'h07;
            16'd25056: data <= 8'hE0;
            16'd25057: data <= 8'h07;
            16'd25058: data <= 8'hE0;
            16'd25059: data <= 8'h07;
            16'd25060: data <= 8'hE0;
            16'd25061: data <= 8'h07;
            16'd25062: data <= 8'hE0;
            16'd25063: data <= 8'h07;
            16'd25064: data <= 8'hE0;
            16'd25065: data <= 8'h07;
            16'd25066: data <= 8'hE0;
            16'd25067: data <= 8'h07;
            16'd25068: data <= 8'hE0;
            16'd25069: data <= 8'h07;
            16'd25070: data <= 8'hE0;
            16'd25071: data <= 8'h07;
            16'd25072: data <= 8'hE0;
            16'd25073: data <= 8'h07;
            16'd25074: data <= 8'hE0;
            16'd25075: data <= 8'h07;
            16'd25076: data <= 8'hE0;
            16'd25077: data <= 8'h07;
            16'd25078: data <= 8'hE0;
            16'd25079: data <= 8'h07;
            16'd25080: data <= 8'hFF;
            16'd25081: data <= 8'hFF;
            16'd25082: data <= 8'hE0;
            16'd25083: data <= 8'h07;
            16'd25084: data <= 8'hE0;
            16'd25085: data <= 8'h07;
            16'd25086: data <= 8'hE0;
            16'd25087: data <= 8'h07;
            16'd25088: data <= 8'hE0;
            16'd25089: data <= 8'h07;
            16'd25090: data <= 8'hE0;
            16'd25091: data <= 8'h07;
            16'd25092: data <= 8'hE0;
            16'd25093: data <= 8'h07;
            16'd25094: data <= 8'hE0;
            16'd25095: data <= 8'h07;
            16'd25096: data <= 8'hE0;
            16'd25097: data <= 8'h07;
            16'd25098: data <= 8'hE0;
            16'd25099: data <= 8'h07;
            16'd25100: data <= 8'hE0;
            16'd25101: data <= 8'h07;
            16'd25102: data <= 8'hE0;
            16'd25103: data <= 8'h07;
            16'd25104: data <= 8'hE0;
            16'd25105: data <= 8'h07;
            16'd25106: data <= 8'hE0;
            16'd25107: data <= 8'h07;
            16'd25108: data <= 8'hE0;
            16'd25109: data <= 8'h07;
            16'd25110: data <= 8'hE0;
            16'd25111: data <= 8'h07;
            16'd25112: data <= 8'hE0;
            16'd25113: data <= 8'h07;
            16'd25114: data <= 8'hE0;
            16'd25115: data <= 8'h07;
            16'd25116: data <= 8'hE0;
            16'd25117: data <= 8'h07;
            16'd25118: data <= 8'hE0;
            16'd25119: data <= 8'h07;
            16'd25120: data <= 8'hFF;
            16'd25121: data <= 8'hFF;
            16'd25122: data <= 8'hE0;
            16'd25123: data <= 8'h07;
            16'd25124: data <= 8'hE0;
            16'd25125: data <= 8'h07;
            16'd25126: data <= 8'hE0;
            16'd25127: data <= 8'h07;
            16'd25128: data <= 8'hE0;
            16'd25129: data <= 8'h07;
            16'd25130: data <= 8'hE0;
            16'd25131: data <= 8'h07;
            16'd25132: data <= 8'hE0;
            16'd25133: data <= 8'h07;
            16'd25134: data <= 8'hE0;
            16'd25135: data <= 8'h07;
            16'd25136: data <= 8'hE0;
            16'd25137: data <= 8'h07;
            16'd25138: data <= 8'hE0;
            16'd25139: data <= 8'h07;
            16'd25140: data <= 8'hE0;
            16'd25141: data <= 8'h07;
            16'd25142: data <= 8'hE0;
            16'd25143: data <= 8'h07;
            16'd25144: data <= 8'hE0;
            16'd25145: data <= 8'h07;
            16'd25146: data <= 8'hE0;
            16'd25147: data <= 8'h07;
            16'd25148: data <= 8'hE0;
            16'd25149: data <= 8'h07;
            16'd25150: data <= 8'hE0;
            16'd25151: data <= 8'h07;
            16'd25152: data <= 8'hE0;
            16'd25153: data <= 8'h07;
            16'd25154: data <= 8'hE0;
            16'd25155: data <= 8'h07;
            16'd25156: data <= 8'hE0;
            16'd25157: data <= 8'h07;
            16'd25158: data <= 8'hE0;
            16'd25159: data <= 8'h07;
            16'd25160: data <= 8'hFF;
            16'd25161: data <= 8'hFF;
            16'd25162: data <= 8'hE0;
            16'd25163: data <= 8'h07;
            16'd25164: data <= 8'hE0;
            16'd25165: data <= 8'h07;
            16'd25166: data <= 8'hE0;
            16'd25167: data <= 8'h07;
            16'd25168: data <= 8'hE0;
            16'd25169: data <= 8'h07;
            16'd25170: data <= 8'hE0;
            16'd25171: data <= 8'h07;
            16'd25172: data <= 8'hE0;
            16'd25173: data <= 8'h07;
            16'd25174: data <= 8'hE0;
            16'd25175: data <= 8'h07;
            16'd25176: data <= 8'hE0;
            16'd25177: data <= 8'h07;
            16'd25178: data <= 8'hE0;
            16'd25179: data <= 8'h07;
            16'd25180: data <= 8'hE0;
            16'd25181: data <= 8'h07;
            16'd25182: data <= 8'hE0;
            16'd25183: data <= 8'h07;
            16'd25184: data <= 8'hE0;
            16'd25185: data <= 8'h07;
            16'd25186: data <= 8'hE0;
            16'd25187: data <= 8'h07;
            16'd25188: data <= 8'hE0;
            16'd25189: data <= 8'h07;
            16'd25190: data <= 8'hE0;
            16'd25191: data <= 8'h07;
            16'd25192: data <= 8'hE0;
            16'd25193: data <= 8'h07;
            16'd25194: data <= 8'hE0;
            16'd25195: data <= 8'h07;
            16'd25196: data <= 8'hE0;
            16'd25197: data <= 8'h07;
            16'd25198: data <= 8'hE0;
            16'd25199: data <= 8'h07;
            16'd25200: data <= 8'hFF;
            16'd25201: data <= 8'hFF;
            16'd25202: data <= 8'hE0;
            16'd25203: data <= 8'h07;
            16'd25204: data <= 8'hE0;
            16'd25205: data <= 8'h07;
            16'd25206: data <= 8'hE0;
            16'd25207: data <= 8'h07;
            16'd25208: data <= 8'hE0;
            16'd25209: data <= 8'h07;
            16'd25210: data <= 8'hE0;
            16'd25211: data <= 8'h07;
            16'd25212: data <= 8'hE0;
            16'd25213: data <= 8'h07;
            16'd25214: data <= 8'hE0;
            16'd25215: data <= 8'h07;
            16'd25216: data <= 8'hE0;
            16'd25217: data <= 8'h07;
            16'd25218: data <= 8'hE0;
            16'd25219: data <= 8'h07;
            16'd25220: data <= 8'hE0;
            16'd25221: data <= 8'h07;
            16'd25222: data <= 8'hE0;
            16'd25223: data <= 8'h07;
            16'd25224: data <= 8'hE0;
            16'd25225: data <= 8'h07;
            16'd25226: data <= 8'hE0;
            16'd25227: data <= 8'h07;
            16'd25228: data <= 8'hE0;
            16'd25229: data <= 8'h07;
            16'd25230: data <= 8'hE0;
            16'd25231: data <= 8'h07;
            16'd25232: data <= 8'hE0;
            16'd25233: data <= 8'h07;
            16'd25234: data <= 8'hE0;
            16'd25235: data <= 8'h07;
            16'd25236: data <= 8'hE0;
            16'd25237: data <= 8'h07;
            16'd25238: data <= 8'hE0;
            16'd25239: data <= 8'h07;
            16'd25240: data <= 8'hFF;
            16'd25241: data <= 8'hFF;
            16'd25242: data <= 8'hE0;
            16'd25243: data <= 8'h07;
            16'd25244: data <= 8'hE0;
            16'd25245: data <= 8'h07;
            16'd25246: data <= 8'hE0;
            16'd25247: data <= 8'h07;
            16'd25248: data <= 8'hE0;
            16'd25249: data <= 8'h07;
            16'd25250: data <= 8'hE0;
            16'd25251: data <= 8'h07;
            16'd25252: data <= 8'hE0;
            16'd25253: data <= 8'h07;
            16'd25254: data <= 8'hE0;
            16'd25255: data <= 8'h07;
            16'd25256: data <= 8'hE0;
            16'd25257: data <= 8'h07;
            16'd25258: data <= 8'hE0;
            16'd25259: data <= 8'h07;
            16'd25260: data <= 8'hE0;
            16'd25261: data <= 8'h07;
            16'd25262: data <= 8'hE0;
            16'd25263: data <= 8'h07;
            16'd25264: data <= 8'hE0;
            16'd25265: data <= 8'h07;
            16'd25266: data <= 8'hE0;
            16'd25267: data <= 8'h07;
            16'd25268: data <= 8'hE0;
            16'd25269: data <= 8'h07;
            16'd25270: data <= 8'hE0;
            16'd25271: data <= 8'h07;
            16'd25272: data <= 8'hE0;
            16'd25273: data <= 8'h07;
            16'd25274: data <= 8'hE0;
            16'd25275: data <= 8'h07;
            16'd25276: data <= 8'hE0;
            16'd25277: data <= 8'h07;
            16'd25278: data <= 8'hE0;
            16'd25279: data <= 8'h07;
            16'd25280: data <= 8'hFF;
            16'd25281: data <= 8'hFF;
            16'd25282: data <= 8'hE0;
            16'd25283: data <= 8'h07;
            16'd25284: data <= 8'hE0;
            16'd25285: data <= 8'h07;
            16'd25286: data <= 8'hE0;
            16'd25287: data <= 8'h07;
            16'd25288: data <= 8'hE0;
            16'd25289: data <= 8'h07;
            16'd25290: data <= 8'hE0;
            16'd25291: data <= 8'h07;
            16'd25292: data <= 8'hE0;
            16'd25293: data <= 8'h07;
            16'd25294: data <= 8'hE0;
            16'd25295: data <= 8'h07;
            16'd25296: data <= 8'hE0;
            16'd25297: data <= 8'h07;
            16'd25298: data <= 8'hE0;
            16'd25299: data <= 8'h07;
            16'd25300: data <= 8'hE0;
            16'd25301: data <= 8'h07;
            16'd25302: data <= 8'hE0;
            16'd25303: data <= 8'h07;
            16'd25304: data <= 8'hE0;
            16'd25305: data <= 8'h07;
            16'd25306: data <= 8'hE0;
            16'd25307: data <= 8'h07;
            16'd25308: data <= 8'hE0;
            16'd25309: data <= 8'h07;
            16'd25310: data <= 8'hE0;
            16'd25311: data <= 8'h07;
            16'd25312: data <= 8'hE0;
            16'd25313: data <= 8'h07;
            16'd25314: data <= 8'hE0;
            16'd25315: data <= 8'h07;
            16'd25316: data <= 8'hE0;
            16'd25317: data <= 8'h07;
            16'd25318: data <= 8'hE0;
            16'd25319: data <= 8'h07;
            16'd25320: data <= 8'hFF;
            16'd25321: data <= 8'hFF;
            16'd25322: data <= 8'hE0;
            16'd25323: data <= 8'h07;
            16'd25324: data <= 8'hE0;
            16'd25325: data <= 8'h07;
            16'd25326: data <= 8'hE0;
            16'd25327: data <= 8'h07;
            16'd25328: data <= 8'hE0;
            16'd25329: data <= 8'h07;
            16'd25330: data <= 8'hE0;
            16'd25331: data <= 8'h07;
            16'd25332: data <= 8'hE0;
            16'd25333: data <= 8'h07;
            16'd25334: data <= 8'hE0;
            16'd25335: data <= 8'h07;
            16'd25336: data <= 8'hE0;
            16'd25337: data <= 8'h07;
            16'd25338: data <= 8'hE0;
            16'd25339: data <= 8'h07;
            16'd25340: data <= 8'hE0;
            16'd25341: data <= 8'h07;
            16'd25342: data <= 8'hE0;
            16'd25343: data <= 8'h07;
            16'd25344: data <= 8'hE0;
            16'd25345: data <= 8'h07;
            16'd25346: data <= 8'hE0;
            16'd25347: data <= 8'h07;
            16'd25348: data <= 8'hE0;
            16'd25349: data <= 8'h07;
            16'd25350: data <= 8'hE0;
            16'd25351: data <= 8'h07;
            16'd25352: data <= 8'hE0;
            16'd25353: data <= 8'h07;
            16'd25354: data <= 8'hE0;
            16'd25355: data <= 8'h07;
            16'd25356: data <= 8'hE0;
            16'd25357: data <= 8'h07;
            16'd25358: data <= 8'hE0;
            16'd25359: data <= 8'h07;
            16'd25360: data <= 8'hFF;
            16'd25361: data <= 8'hFF;
            16'd25362: data <= 8'hE0;
            16'd25363: data <= 8'h07;
            16'd25364: data <= 8'hE0;
            16'd25365: data <= 8'h07;
            16'd25366: data <= 8'hE0;
            16'd25367: data <= 8'h07;
            16'd25368: data <= 8'hE0;
            16'd25369: data <= 8'h07;
            16'd25370: data <= 8'hE0;
            16'd25371: data <= 8'h07;
            16'd25372: data <= 8'hE0;
            16'd25373: data <= 8'h07;
            16'd25374: data <= 8'hE0;
            16'd25375: data <= 8'h07;
            16'd25376: data <= 8'hE0;
            16'd25377: data <= 8'h07;
            16'd25378: data <= 8'hE0;
            16'd25379: data <= 8'h07;
            16'd25380: data <= 8'hE0;
            16'd25381: data <= 8'h07;
            16'd25382: data <= 8'hE0;
            16'd25383: data <= 8'h07;
            16'd25384: data <= 8'hE0;
            16'd25385: data <= 8'h07;
            16'd25386: data <= 8'hE0;
            16'd25387: data <= 8'h07;
            16'd25388: data <= 8'hE0;
            16'd25389: data <= 8'h07;
            16'd25390: data <= 8'hE0;
            16'd25391: data <= 8'h07;
            16'd25392: data <= 8'hE0;
            16'd25393: data <= 8'h07;
            16'd25394: data <= 8'hE0;
            16'd25395: data <= 8'h07;
            16'd25396: data <= 8'hE0;
            16'd25397: data <= 8'h07;
            16'd25398: data <= 8'hE0;
            16'd25399: data <= 8'h07;
            16'd25400: data <= 8'hFF;
            16'd25401: data <= 8'hFF;
            16'd25402: data <= 8'hE0;
            16'd25403: data <= 8'h07;
            16'd25404: data <= 8'hE0;
            16'd25405: data <= 8'h07;
            16'd25406: data <= 8'hE0;
            16'd25407: data <= 8'h07;
            16'd25408: data <= 8'hE0;
            16'd25409: data <= 8'h07;
            16'd25410: data <= 8'hE0;
            16'd25411: data <= 8'h07;
            16'd25412: data <= 8'hE0;
            16'd25413: data <= 8'h07;
            16'd25414: data <= 8'hE0;
            16'd25415: data <= 8'h07;
            16'd25416: data <= 8'hE0;
            16'd25417: data <= 8'h07;
            16'd25418: data <= 8'hE0;
            16'd25419: data <= 8'h07;
            16'd25420: data <= 8'hE0;
            16'd25421: data <= 8'h07;
            16'd25422: data <= 8'hE0;
            16'd25423: data <= 8'h07;
            16'd25424: data <= 8'hE0;
            16'd25425: data <= 8'h07;
            16'd25426: data <= 8'hE0;
            16'd25427: data <= 8'h07;
            16'd25428: data <= 8'hE0;
            16'd25429: data <= 8'h07;
            16'd25430: data <= 8'hE0;
            16'd25431: data <= 8'h07;
            16'd25432: data <= 8'hE0;
            16'd25433: data <= 8'h07;
            16'd25434: data <= 8'hE0;
            16'd25435: data <= 8'h07;
            16'd25436: data <= 8'hE0;
            16'd25437: data <= 8'h07;
            16'd25438: data <= 8'hE0;
            16'd25439: data <= 8'h07;
            16'd25440: data <= 8'hFF;
            16'd25441: data <= 8'hFF;
            16'd25442: data <= 8'h1F;
            16'd25443: data <= 8'h00;
            16'd25444: data <= 8'h1F;
            16'd25445: data <= 8'h00;
            16'd25446: data <= 8'h1F;
            16'd25447: data <= 8'h00;
            16'd25448: data <= 8'h1F;
            16'd25449: data <= 8'h00;
            16'd25450: data <= 8'h1F;
            16'd25451: data <= 8'h00;
            16'd25452: data <= 8'h1F;
            16'd25453: data <= 8'h00;
            16'd25454: data <= 8'h1F;
            16'd25455: data <= 8'h00;
            16'd25456: data <= 8'h1F;
            16'd25457: data <= 8'h00;
            16'd25458: data <= 8'h1F;
            16'd25459: data <= 8'h00;
            16'd25460: data <= 8'h1F;
            16'd25461: data <= 8'h00;
            16'd25462: data <= 8'h1F;
            16'd25463: data <= 8'h00;
            16'd25464: data <= 8'h1F;
            16'd25465: data <= 8'h00;
            16'd25466: data <= 8'h1F;
            16'd25467: data <= 8'h00;
            16'd25468: data <= 8'h1F;
            16'd25469: data <= 8'h00;
            16'd25470: data <= 8'h1F;
            16'd25471: data <= 8'h00;
            16'd25472: data <= 8'h1F;
            16'd25473: data <= 8'h00;
            16'd25474: data <= 8'h1F;
            16'd25475: data <= 8'h00;
            16'd25476: data <= 8'h1F;
            16'd25477: data <= 8'h00;
            16'd25478: data <= 8'h1F;
            16'd25479: data <= 8'h00;
            16'd25480: data <= 8'hFF;
            16'd25481: data <= 8'hFF;
            16'd25482: data <= 8'h1F;
            16'd25483: data <= 8'h00;
            16'd25484: data <= 8'h1F;
            16'd25485: data <= 8'h00;
            16'd25486: data <= 8'h1F;
            16'd25487: data <= 8'h00;
            16'd25488: data <= 8'h1F;
            16'd25489: data <= 8'h00;
            16'd25490: data <= 8'h1F;
            16'd25491: data <= 8'h00;
            16'd25492: data <= 8'h1F;
            16'd25493: data <= 8'h00;
            16'd25494: data <= 8'h1F;
            16'd25495: data <= 8'h00;
            16'd25496: data <= 8'h1F;
            16'd25497: data <= 8'h00;
            16'd25498: data <= 8'h1F;
            16'd25499: data <= 8'h00;
            16'd25500: data <= 8'h1F;
            16'd25501: data <= 8'h00;
            16'd25502: data <= 8'h1F;
            16'd25503: data <= 8'h00;
            16'd25504: data <= 8'h1F;
            16'd25505: data <= 8'h00;
            16'd25506: data <= 8'h1F;
            16'd25507: data <= 8'h00;
            16'd25508: data <= 8'h1F;
            16'd25509: data <= 8'h00;
            16'd25510: data <= 8'h1F;
            16'd25511: data <= 8'h00;
            16'd25512: data <= 8'h1F;
            16'd25513: data <= 8'h00;
            16'd25514: data <= 8'h1F;
            16'd25515: data <= 8'h00;
            16'd25516: data <= 8'h1F;
            16'd25517: data <= 8'h00;
            16'd25518: data <= 8'h1F;
            16'd25519: data <= 8'h00;
            16'd25520: data <= 8'hFF;
            16'd25521: data <= 8'hFF;
            16'd25522: data <= 8'h1F;
            16'd25523: data <= 8'h00;
            16'd25524: data <= 8'h1F;
            16'd25525: data <= 8'h00;
            16'd25526: data <= 8'h1F;
            16'd25527: data <= 8'h00;
            16'd25528: data <= 8'h1F;
            16'd25529: data <= 8'h00;
            16'd25530: data <= 8'h1F;
            16'd25531: data <= 8'h00;
            16'd25532: data <= 8'h1F;
            16'd25533: data <= 8'h00;
            16'd25534: data <= 8'h1F;
            16'd25535: data <= 8'h00;
            16'd25536: data <= 8'h1F;
            16'd25537: data <= 8'h00;
            16'd25538: data <= 8'h1F;
            16'd25539: data <= 8'h00;
            16'd25540: data <= 8'h1F;
            16'd25541: data <= 8'h00;
            16'd25542: data <= 8'h1F;
            16'd25543: data <= 8'h00;
            16'd25544: data <= 8'h1F;
            16'd25545: data <= 8'h00;
            16'd25546: data <= 8'h1F;
            16'd25547: data <= 8'h00;
            16'd25548: data <= 8'h1F;
            16'd25549: data <= 8'h00;
            16'd25550: data <= 8'h1F;
            16'd25551: data <= 8'h00;
            16'd25552: data <= 8'h1F;
            16'd25553: data <= 8'h00;
            16'd25554: data <= 8'h1F;
            16'd25555: data <= 8'h00;
            16'd25556: data <= 8'h1F;
            16'd25557: data <= 8'h00;
            16'd25558: data <= 8'h1F;
            16'd25559: data <= 8'h00;
            16'd25560: data <= 8'hFF;
            16'd25561: data <= 8'hFF;
            16'd25562: data <= 8'h1F;
            16'd25563: data <= 8'h00;
            16'd25564: data <= 8'h1F;
            16'd25565: data <= 8'h00;
            16'd25566: data <= 8'h1F;
            16'd25567: data <= 8'h00;
            16'd25568: data <= 8'h1F;
            16'd25569: data <= 8'h00;
            16'd25570: data <= 8'h1F;
            16'd25571: data <= 8'h00;
            16'd25572: data <= 8'h1F;
            16'd25573: data <= 8'h00;
            16'd25574: data <= 8'h1F;
            16'd25575: data <= 8'h00;
            16'd25576: data <= 8'h1F;
            16'd25577: data <= 8'h00;
            16'd25578: data <= 8'h1F;
            16'd25579: data <= 8'h00;
            16'd25580: data <= 8'h1F;
            16'd25581: data <= 8'h00;
            16'd25582: data <= 8'h1F;
            16'd25583: data <= 8'h00;
            16'd25584: data <= 8'h1F;
            16'd25585: data <= 8'h00;
            16'd25586: data <= 8'h1F;
            16'd25587: data <= 8'h00;
            16'd25588: data <= 8'h1F;
            16'd25589: data <= 8'h00;
            16'd25590: data <= 8'h1F;
            16'd25591: data <= 8'h00;
            16'd25592: data <= 8'h1F;
            16'd25593: data <= 8'h00;
            16'd25594: data <= 8'h1F;
            16'd25595: data <= 8'h00;
            16'd25596: data <= 8'h1F;
            16'd25597: data <= 8'h00;
            16'd25598: data <= 8'h1F;
            16'd25599: data <= 8'h00;
            16'd25600: data <= 8'hFF;
            16'd25601: data <= 8'hFF;
            16'd25602: data <= 8'h1F;
            16'd25603: data <= 8'h00;
            16'd25604: data <= 8'h1F;
            16'd25605: data <= 8'h00;
            16'd25606: data <= 8'h1F;
            16'd25607: data <= 8'h00;
            16'd25608: data <= 8'h1F;
            16'd25609: data <= 8'h00;
            16'd25610: data <= 8'h1F;
            16'd25611: data <= 8'h00;
            16'd25612: data <= 8'h1F;
            16'd25613: data <= 8'h00;
            16'd25614: data <= 8'h1F;
            16'd25615: data <= 8'h00;
            16'd25616: data <= 8'h1F;
            16'd25617: data <= 8'h00;
            16'd25618: data <= 8'h1F;
            16'd25619: data <= 8'h00;
            16'd25620: data <= 8'h1F;
            16'd25621: data <= 8'h00;
            16'd25622: data <= 8'h1F;
            16'd25623: data <= 8'h00;
            16'd25624: data <= 8'h1F;
            16'd25625: data <= 8'h00;
            16'd25626: data <= 8'h1F;
            16'd25627: data <= 8'h00;
            16'd25628: data <= 8'h1F;
            16'd25629: data <= 8'h00;
            16'd25630: data <= 8'h1F;
            16'd25631: data <= 8'h00;
            16'd25632: data <= 8'h1F;
            16'd25633: data <= 8'h00;
            16'd25634: data <= 8'h1F;
            16'd25635: data <= 8'h00;
            16'd25636: data <= 8'h1F;
            16'd25637: data <= 8'h00;
            16'd25638: data <= 8'h1F;
            16'd25639: data <= 8'h00;
            16'd25640: data <= 8'hFF;
            16'd25641: data <= 8'hFF;
            16'd25642: data <= 8'h1F;
            16'd25643: data <= 8'h00;
            16'd25644: data <= 8'h1F;
            16'd25645: data <= 8'h00;
            16'd25646: data <= 8'h1F;
            16'd25647: data <= 8'h00;
            16'd25648: data <= 8'h1F;
            16'd25649: data <= 8'h00;
            16'd25650: data <= 8'h1F;
            16'd25651: data <= 8'h00;
            16'd25652: data <= 8'h1F;
            16'd25653: data <= 8'h00;
            16'd25654: data <= 8'h1F;
            16'd25655: data <= 8'h00;
            16'd25656: data <= 8'h1F;
            16'd25657: data <= 8'h00;
            16'd25658: data <= 8'h1F;
            16'd25659: data <= 8'h00;
            16'd25660: data <= 8'h1F;
            16'd25661: data <= 8'h00;
            16'd25662: data <= 8'h1F;
            16'd25663: data <= 8'h00;
            16'd25664: data <= 8'h1F;
            16'd25665: data <= 8'h00;
            16'd25666: data <= 8'h1F;
            16'd25667: data <= 8'h00;
            16'd25668: data <= 8'h1F;
            16'd25669: data <= 8'h00;
            16'd25670: data <= 8'h1F;
            16'd25671: data <= 8'h00;
            16'd25672: data <= 8'h1F;
            16'd25673: data <= 8'h00;
            16'd25674: data <= 8'h1F;
            16'd25675: data <= 8'h00;
            16'd25676: data <= 8'h1F;
            16'd25677: data <= 8'h00;
            16'd25678: data <= 8'h1F;
            16'd25679: data <= 8'h00;
            16'd25680: data <= 8'hFF;
            16'd25681: data <= 8'hFF;
            16'd25682: data <= 8'h1F;
            16'd25683: data <= 8'h00;
            16'd25684: data <= 8'h1F;
            16'd25685: data <= 8'h00;
            16'd25686: data <= 8'h1F;
            16'd25687: data <= 8'h00;
            16'd25688: data <= 8'h1F;
            16'd25689: data <= 8'h00;
            16'd25690: data <= 8'h1F;
            16'd25691: data <= 8'h00;
            16'd25692: data <= 8'h1F;
            16'd25693: data <= 8'h00;
            16'd25694: data <= 8'h1F;
            16'd25695: data <= 8'h00;
            16'd25696: data <= 8'h1F;
            16'd25697: data <= 8'h00;
            16'd25698: data <= 8'h1F;
            16'd25699: data <= 8'h00;
            16'd25700: data <= 8'h1F;
            16'd25701: data <= 8'h00;
            16'd25702: data <= 8'h1F;
            16'd25703: data <= 8'h00;
            16'd25704: data <= 8'h1F;
            16'd25705: data <= 8'h00;
            16'd25706: data <= 8'h1F;
            16'd25707: data <= 8'h00;
            16'd25708: data <= 8'h1F;
            16'd25709: data <= 8'h00;
            16'd25710: data <= 8'h1F;
            16'd25711: data <= 8'h00;
            16'd25712: data <= 8'h1F;
            16'd25713: data <= 8'h00;
            16'd25714: data <= 8'h1F;
            16'd25715: data <= 8'h00;
            16'd25716: data <= 8'h1F;
            16'd25717: data <= 8'h00;
            16'd25718: data <= 8'h1F;
            16'd25719: data <= 8'h00;
            16'd25720: data <= 8'hFF;
            16'd25721: data <= 8'hFF;
            16'd25722: data <= 8'h1F;
            16'd25723: data <= 8'h00;
            16'd25724: data <= 8'h1F;
            16'd25725: data <= 8'h00;
            16'd25726: data <= 8'h1F;
            16'd25727: data <= 8'h00;
            16'd25728: data <= 8'h1F;
            16'd25729: data <= 8'h00;
            16'd25730: data <= 8'h1F;
            16'd25731: data <= 8'h00;
            16'd25732: data <= 8'h1F;
            16'd25733: data <= 8'h00;
            16'd25734: data <= 8'h1F;
            16'd25735: data <= 8'h00;
            16'd25736: data <= 8'h1F;
            16'd25737: data <= 8'h00;
            16'd25738: data <= 8'h1F;
            16'd25739: data <= 8'h00;
            16'd25740: data <= 8'h1F;
            16'd25741: data <= 8'h00;
            16'd25742: data <= 8'h1F;
            16'd25743: data <= 8'h00;
            16'd25744: data <= 8'h1F;
            16'd25745: data <= 8'h00;
            16'd25746: data <= 8'h1F;
            16'd25747: data <= 8'h00;
            16'd25748: data <= 8'h1F;
            16'd25749: data <= 8'h00;
            16'd25750: data <= 8'h1F;
            16'd25751: data <= 8'h00;
            16'd25752: data <= 8'h1F;
            16'd25753: data <= 8'h00;
            16'd25754: data <= 8'h1F;
            16'd25755: data <= 8'h00;
            16'd25756: data <= 8'h1F;
            16'd25757: data <= 8'h00;
            16'd25758: data <= 8'h1F;
            16'd25759: data <= 8'h00;
            16'd25760: data <= 8'hFF;
            16'd25761: data <= 8'hFF;
            16'd25762: data <= 8'h1F;
            16'd25763: data <= 8'h00;
            16'd25764: data <= 8'h1F;
            16'd25765: data <= 8'h00;
            16'd25766: data <= 8'h1F;
            16'd25767: data <= 8'h00;
            16'd25768: data <= 8'h1F;
            16'd25769: data <= 8'h00;
            16'd25770: data <= 8'h1F;
            16'd25771: data <= 8'h00;
            16'd25772: data <= 8'h1F;
            16'd25773: data <= 8'h00;
            16'd25774: data <= 8'h1F;
            16'd25775: data <= 8'h00;
            16'd25776: data <= 8'h1F;
            16'd25777: data <= 8'h00;
            16'd25778: data <= 8'h1F;
            16'd25779: data <= 8'h00;
            16'd25780: data <= 8'h1F;
            16'd25781: data <= 8'h00;
            16'd25782: data <= 8'h1F;
            16'd25783: data <= 8'h00;
            16'd25784: data <= 8'h1F;
            16'd25785: data <= 8'h00;
            16'd25786: data <= 8'h1F;
            16'd25787: data <= 8'h00;
            16'd25788: data <= 8'h1F;
            16'd25789: data <= 8'h00;
            16'd25790: data <= 8'h1F;
            16'd25791: data <= 8'h00;
            16'd25792: data <= 8'h1F;
            16'd25793: data <= 8'h00;
            16'd25794: data <= 8'h1F;
            16'd25795: data <= 8'h00;
            16'd25796: data <= 8'h1F;
            16'd25797: data <= 8'h00;
            16'd25798: data <= 8'h1F;
            16'd25799: data <= 8'h00;
            16'd25800: data <= 8'hFF;
            16'd25801: data <= 8'hFF;
            16'd25802: data <= 8'h1F;
            16'd25803: data <= 8'h00;
            16'd25804: data <= 8'h1F;
            16'd25805: data <= 8'h00;
            16'd25806: data <= 8'h1F;
            16'd25807: data <= 8'h00;
            16'd25808: data <= 8'h1F;
            16'd25809: data <= 8'h00;
            16'd25810: data <= 8'h1F;
            16'd25811: data <= 8'h00;
            16'd25812: data <= 8'h1F;
            16'd25813: data <= 8'h00;
            16'd25814: data <= 8'h1F;
            16'd25815: data <= 8'h00;
            16'd25816: data <= 8'h1F;
            16'd25817: data <= 8'h00;
            16'd25818: data <= 8'h1F;
            16'd25819: data <= 8'h00;
            16'd25820: data <= 8'h1F;
            16'd25821: data <= 8'h00;
            16'd25822: data <= 8'h1F;
            16'd25823: data <= 8'h00;
            16'd25824: data <= 8'h1F;
            16'd25825: data <= 8'h00;
            16'd25826: data <= 8'h1F;
            16'd25827: data <= 8'h00;
            16'd25828: data <= 8'h1F;
            16'd25829: data <= 8'h00;
            16'd25830: data <= 8'h1F;
            16'd25831: data <= 8'h00;
            16'd25832: data <= 8'h1F;
            16'd25833: data <= 8'h00;
            16'd25834: data <= 8'h1F;
            16'd25835: data <= 8'h00;
            16'd25836: data <= 8'h1F;
            16'd25837: data <= 8'h00;
            16'd25838: data <= 8'h1F;
            16'd25839: data <= 8'h00;
            16'd25840: data <= 8'hFF;
            16'd25841: data <= 8'hFF;
            16'd25842: data <= 8'h1F;
            16'd25843: data <= 8'h00;
            16'd25844: data <= 8'h1F;
            16'd25845: data <= 8'h00;
            16'd25846: data <= 8'h1F;
            16'd25847: data <= 8'h00;
            16'd25848: data <= 8'h1F;
            16'd25849: data <= 8'h00;
            16'd25850: data <= 8'h1F;
            16'd25851: data <= 8'h00;
            16'd25852: data <= 8'h1F;
            16'd25853: data <= 8'h00;
            16'd25854: data <= 8'h1F;
            16'd25855: data <= 8'h00;
            16'd25856: data <= 8'h1F;
            16'd25857: data <= 8'h00;
            16'd25858: data <= 8'h1F;
            16'd25859: data <= 8'h00;
            16'd25860: data <= 8'h1F;
            16'd25861: data <= 8'h00;
            16'd25862: data <= 8'h1F;
            16'd25863: data <= 8'h00;
            16'd25864: data <= 8'h1F;
            16'd25865: data <= 8'h00;
            16'd25866: data <= 8'h1F;
            16'd25867: data <= 8'h00;
            16'd25868: data <= 8'h1F;
            16'd25869: data <= 8'h00;
            16'd25870: data <= 8'h1F;
            16'd25871: data <= 8'h00;
            16'd25872: data <= 8'h1F;
            16'd25873: data <= 8'h00;
            16'd25874: data <= 8'h1F;
            16'd25875: data <= 8'h00;
            16'd25876: data <= 8'h1F;
            16'd25877: data <= 8'h00;
            16'd25878: data <= 8'h1F;
            16'd25879: data <= 8'h00;
            16'd25880: data <= 8'hFF;
            16'd25881: data <= 8'hFF;
            16'd25882: data <= 8'h1F;
            16'd25883: data <= 8'h00;
            16'd25884: data <= 8'h1F;
            16'd25885: data <= 8'h00;
            16'd25886: data <= 8'h1F;
            16'd25887: data <= 8'h00;
            16'd25888: data <= 8'h1F;
            16'd25889: data <= 8'h00;
            16'd25890: data <= 8'h1F;
            16'd25891: data <= 8'h00;
            16'd25892: data <= 8'h1F;
            16'd25893: data <= 8'h00;
            16'd25894: data <= 8'h1F;
            16'd25895: data <= 8'h00;
            16'd25896: data <= 8'h1F;
            16'd25897: data <= 8'h00;
            16'd25898: data <= 8'h1F;
            16'd25899: data <= 8'h00;
            16'd25900: data <= 8'h1F;
            16'd25901: data <= 8'h00;
            16'd25902: data <= 8'h1F;
            16'd25903: data <= 8'h00;
            16'd25904: data <= 8'h1F;
            16'd25905: data <= 8'h00;
            16'd25906: data <= 8'h1F;
            16'd25907: data <= 8'h00;
            16'd25908: data <= 8'h1F;
            16'd25909: data <= 8'h00;
            16'd25910: data <= 8'h1F;
            16'd25911: data <= 8'h00;
            16'd25912: data <= 8'h1F;
            16'd25913: data <= 8'h00;
            16'd25914: data <= 8'h1F;
            16'd25915: data <= 8'h00;
            16'd25916: data <= 8'h1F;
            16'd25917: data <= 8'h00;
            16'd25918: data <= 8'h1F;
            16'd25919: data <= 8'h00;
            16'd25920: data <= 8'hFF;
            16'd25921: data <= 8'hFF;
            16'd25922: data <= 8'h1F;
            16'd25923: data <= 8'h00;
            16'd25924: data <= 8'h1F;
            16'd25925: data <= 8'h00;
            16'd25926: data <= 8'h1F;
            16'd25927: data <= 8'h00;
            16'd25928: data <= 8'h1F;
            16'd25929: data <= 8'h00;
            16'd25930: data <= 8'h1F;
            16'd25931: data <= 8'h00;
            16'd25932: data <= 8'h1F;
            16'd25933: data <= 8'h00;
            16'd25934: data <= 8'h1F;
            16'd25935: data <= 8'h00;
            16'd25936: data <= 8'h1F;
            16'd25937: data <= 8'h00;
            16'd25938: data <= 8'h1F;
            16'd25939: data <= 8'h00;
            16'd25940: data <= 8'h1F;
            16'd25941: data <= 8'h00;
            16'd25942: data <= 8'h1F;
            16'd25943: data <= 8'h00;
            16'd25944: data <= 8'h1F;
            16'd25945: data <= 8'h00;
            16'd25946: data <= 8'h1F;
            16'd25947: data <= 8'h00;
            16'd25948: data <= 8'h1F;
            16'd25949: data <= 8'h00;
            16'd25950: data <= 8'h1F;
            16'd25951: data <= 8'h00;
            16'd25952: data <= 8'h1F;
            16'd25953: data <= 8'h00;
            16'd25954: data <= 8'h1F;
            16'd25955: data <= 8'h00;
            16'd25956: data <= 8'h1F;
            16'd25957: data <= 8'h00;
            16'd25958: data <= 8'h1F;
            16'd25959: data <= 8'h00;
            16'd25960: data <= 8'hFF;
            16'd25961: data <= 8'hFF;
            16'd25962: data <= 8'h1F;
            16'd25963: data <= 8'h00;
            16'd25964: data <= 8'h1F;
            16'd25965: data <= 8'h00;
            16'd25966: data <= 8'h1F;
            16'd25967: data <= 8'h00;
            16'd25968: data <= 8'h1F;
            16'd25969: data <= 8'h00;
            16'd25970: data <= 8'h1F;
            16'd25971: data <= 8'h00;
            16'd25972: data <= 8'h1F;
            16'd25973: data <= 8'h00;
            16'd25974: data <= 8'h1F;
            16'd25975: data <= 8'h00;
            16'd25976: data <= 8'h1F;
            16'd25977: data <= 8'h00;
            16'd25978: data <= 8'h1F;
            16'd25979: data <= 8'h00;
            16'd25980: data <= 8'h1F;
            16'd25981: data <= 8'h00;
            16'd25982: data <= 8'h1F;
            16'd25983: data <= 8'h00;
            16'd25984: data <= 8'h1F;
            16'd25985: data <= 8'h00;
            16'd25986: data <= 8'h1F;
            16'd25987: data <= 8'h00;
            16'd25988: data <= 8'h1F;
            16'd25989: data <= 8'h00;
            16'd25990: data <= 8'h1F;
            16'd25991: data <= 8'h00;
            16'd25992: data <= 8'h1F;
            16'd25993: data <= 8'h00;
            16'd25994: data <= 8'h1F;
            16'd25995: data <= 8'h00;
            16'd25996: data <= 8'h1F;
            16'd25997: data <= 8'h00;
            16'd25998: data <= 8'h1F;
            16'd25999: data <= 8'h00;
            16'd26000: data <= 8'hFF;
            16'd26001: data <= 8'hFF;
            16'd26002: data <= 8'h1F;
            16'd26003: data <= 8'h00;
            16'd26004: data <= 8'h1F;
            16'd26005: data <= 8'h00;
            16'd26006: data <= 8'h1F;
            16'd26007: data <= 8'h00;
            16'd26008: data <= 8'h1F;
            16'd26009: data <= 8'h00;
            16'd26010: data <= 8'h1F;
            16'd26011: data <= 8'h00;
            16'd26012: data <= 8'h1F;
            16'd26013: data <= 8'h00;
            16'd26014: data <= 8'h1F;
            16'd26015: data <= 8'h00;
            16'd26016: data <= 8'h1F;
            16'd26017: data <= 8'h00;
            16'd26018: data <= 8'h1F;
            16'd26019: data <= 8'h00;
            16'd26020: data <= 8'h1F;
            16'd26021: data <= 8'h00;
            16'd26022: data <= 8'h1F;
            16'd26023: data <= 8'h00;
            16'd26024: data <= 8'h1F;
            16'd26025: data <= 8'h00;
            16'd26026: data <= 8'h1F;
            16'd26027: data <= 8'h00;
            16'd26028: data <= 8'h1F;
            16'd26029: data <= 8'h00;
            16'd26030: data <= 8'h1F;
            16'd26031: data <= 8'h00;
            16'd26032: data <= 8'h1F;
            16'd26033: data <= 8'h00;
            16'd26034: data <= 8'h1F;
            16'd26035: data <= 8'h00;
            16'd26036: data <= 8'h1F;
            16'd26037: data <= 8'h00;
            16'd26038: data <= 8'h1F;
            16'd26039: data <= 8'h00;
            16'd26040: data <= 8'hFF;
            16'd26041: data <= 8'hFF;
            16'd26042: data <= 8'h1F;
            16'd26043: data <= 8'h00;
            16'd26044: data <= 8'h1F;
            16'd26045: data <= 8'h00;
            16'd26046: data <= 8'h1F;
            16'd26047: data <= 8'h00;
            16'd26048: data <= 8'h1F;
            16'd26049: data <= 8'h00;
            16'd26050: data <= 8'h1F;
            16'd26051: data <= 8'h00;
            16'd26052: data <= 8'h1F;
            16'd26053: data <= 8'h00;
            16'd26054: data <= 8'h1F;
            16'd26055: data <= 8'h00;
            16'd26056: data <= 8'h1F;
            16'd26057: data <= 8'h00;
            16'd26058: data <= 8'h1F;
            16'd26059: data <= 8'h00;
            16'd26060: data <= 8'h1F;
            16'd26061: data <= 8'h00;
            16'd26062: data <= 8'h1F;
            16'd26063: data <= 8'h00;
            16'd26064: data <= 8'h1F;
            16'd26065: data <= 8'h00;
            16'd26066: data <= 8'h1F;
            16'd26067: data <= 8'h00;
            16'd26068: data <= 8'h1F;
            16'd26069: data <= 8'h00;
            16'd26070: data <= 8'h1F;
            16'd26071: data <= 8'h00;
            16'd26072: data <= 8'h1F;
            16'd26073: data <= 8'h00;
            16'd26074: data <= 8'h1F;
            16'd26075: data <= 8'h00;
            16'd26076: data <= 8'h1F;
            16'd26077: data <= 8'h00;
            16'd26078: data <= 8'h1F;
            16'd26079: data <= 8'h00;
            16'd26080: data <= 8'hFF;
            16'd26081: data <= 8'hFF;
            16'd26082: data <= 8'h1F;
            16'd26083: data <= 8'h00;
            16'd26084: data <= 8'h1F;
            16'd26085: data <= 8'h00;
            16'd26086: data <= 8'h1F;
            16'd26087: data <= 8'h00;
            16'd26088: data <= 8'h1F;
            16'd26089: data <= 8'h00;
            16'd26090: data <= 8'h1F;
            16'd26091: data <= 8'h00;
            16'd26092: data <= 8'h1F;
            16'd26093: data <= 8'h00;
            16'd26094: data <= 8'h1F;
            16'd26095: data <= 8'h00;
            16'd26096: data <= 8'h1F;
            16'd26097: data <= 8'h00;
            16'd26098: data <= 8'h1F;
            16'd26099: data <= 8'h00;
            16'd26100: data <= 8'h1F;
            16'd26101: data <= 8'h00;
            16'd26102: data <= 8'h1F;
            16'd26103: data <= 8'h00;
            16'd26104: data <= 8'h1F;
            16'd26105: data <= 8'h00;
            16'd26106: data <= 8'h1F;
            16'd26107: data <= 8'h00;
            16'd26108: data <= 8'h1F;
            16'd26109: data <= 8'h00;
            16'd26110: data <= 8'h1F;
            16'd26111: data <= 8'h00;
            16'd26112: data <= 8'h1F;
            16'd26113: data <= 8'h00;
            16'd26114: data <= 8'h1F;
            16'd26115: data <= 8'h00;
            16'd26116: data <= 8'h1F;
            16'd26117: data <= 8'h00;
            16'd26118: data <= 8'h1F;
            16'd26119: data <= 8'h00;
            16'd26120: data <= 8'hFF;
            16'd26121: data <= 8'hFF;
            16'd26122: data <= 8'h1F;
            16'd26123: data <= 8'h00;
            16'd26124: data <= 8'h1F;
            16'd26125: data <= 8'h00;
            16'd26126: data <= 8'h1F;
            16'd26127: data <= 8'h00;
            16'd26128: data <= 8'h1F;
            16'd26129: data <= 8'h00;
            16'd26130: data <= 8'h1F;
            16'd26131: data <= 8'h00;
            16'd26132: data <= 8'h1F;
            16'd26133: data <= 8'h00;
            16'd26134: data <= 8'h1F;
            16'd26135: data <= 8'h00;
            16'd26136: data <= 8'h1F;
            16'd26137: data <= 8'h00;
            16'd26138: data <= 8'h1F;
            16'd26139: data <= 8'h00;
            16'd26140: data <= 8'h1F;
            16'd26141: data <= 8'h00;
            16'd26142: data <= 8'h1F;
            16'd26143: data <= 8'h00;
            16'd26144: data <= 8'h1F;
            16'd26145: data <= 8'h00;
            16'd26146: data <= 8'h1F;
            16'd26147: data <= 8'h00;
            16'd26148: data <= 8'h1F;
            16'd26149: data <= 8'h00;
            16'd26150: data <= 8'h1F;
            16'd26151: data <= 8'h00;
            16'd26152: data <= 8'h1F;
            16'd26153: data <= 8'h00;
            16'd26154: data <= 8'h1F;
            16'd26155: data <= 8'h00;
            16'd26156: data <= 8'h1F;
            16'd26157: data <= 8'h00;
            16'd26158: data <= 8'h1F;
            16'd26159: data <= 8'h00;
            16'd26160: data <= 8'hFF;
            16'd26161: data <= 8'hFF;
            16'd26162: data <= 8'h1F;
            16'd26163: data <= 8'h00;
            16'd26164: data <= 8'h1F;
            16'd26165: data <= 8'h00;
            16'd26166: data <= 8'h1F;
            16'd26167: data <= 8'h00;
            16'd26168: data <= 8'h1F;
            16'd26169: data <= 8'h00;
            16'd26170: data <= 8'h1F;
            16'd26171: data <= 8'h00;
            16'd26172: data <= 8'h1F;
            16'd26173: data <= 8'h00;
            16'd26174: data <= 8'h1F;
            16'd26175: data <= 8'h00;
            16'd26176: data <= 8'h1F;
            16'd26177: data <= 8'h00;
            16'd26178: data <= 8'h1F;
            16'd26179: data <= 8'h00;
            16'd26180: data <= 8'h1F;
            16'd26181: data <= 8'h00;
            16'd26182: data <= 8'h1F;
            16'd26183: data <= 8'h00;
            16'd26184: data <= 8'h1F;
            16'd26185: data <= 8'h00;
            16'd26186: data <= 8'h1F;
            16'd26187: data <= 8'h00;
            16'd26188: data <= 8'h1F;
            16'd26189: data <= 8'h00;
            16'd26190: data <= 8'h1F;
            16'd26191: data <= 8'h00;
            16'd26192: data <= 8'h1F;
            16'd26193: data <= 8'h00;
            16'd26194: data <= 8'h1F;
            16'd26195: data <= 8'h00;
            16'd26196: data <= 8'h1F;
            16'd26197: data <= 8'h00;
            16'd26198: data <= 8'h1F;
            16'd26199: data <= 8'h00;
            16'd26200: data <= 8'hFF;
            16'd26201: data <= 8'hFF;
            16'd26202: data <= 8'h1F;
            16'd26203: data <= 8'h00;
            16'd26204: data <= 8'h1F;
            16'd26205: data <= 8'h00;
            16'd26206: data <= 8'h1F;
            16'd26207: data <= 8'h00;
            16'd26208: data <= 8'h1F;
            16'd26209: data <= 8'h00;
            16'd26210: data <= 8'h1F;
            16'd26211: data <= 8'h00;
            16'd26212: data <= 8'h1F;
            16'd26213: data <= 8'h00;
            16'd26214: data <= 8'h1F;
            16'd26215: data <= 8'h00;
            16'd26216: data <= 8'h1F;
            16'd26217: data <= 8'h00;
            16'd26218: data <= 8'h1F;
            16'd26219: data <= 8'h00;
            16'd26220: data <= 8'h1F;
            16'd26221: data <= 8'h00;
            16'd26222: data <= 8'h1F;
            16'd26223: data <= 8'h00;
            16'd26224: data <= 8'h1F;
            16'd26225: data <= 8'h00;
            16'd26226: data <= 8'h1F;
            16'd26227: data <= 8'h00;
            16'd26228: data <= 8'h1F;
            16'd26229: data <= 8'h00;
            16'd26230: data <= 8'h1F;
            16'd26231: data <= 8'h00;
            16'd26232: data <= 8'h1F;
            16'd26233: data <= 8'h00;
            16'd26234: data <= 8'h1F;
            16'd26235: data <= 8'h00;
            16'd26236: data <= 8'h1F;
            16'd26237: data <= 8'h00;
            16'd26238: data <= 8'h1F;
            16'd26239: data <= 8'h00;
            16'd26240: data <= 8'hFF;
            16'd26241: data <= 8'hFF;
            16'd26242: data <= 8'h1F;
            16'd26243: data <= 8'h00;
            16'd26244: data <= 8'h1F;
            16'd26245: data <= 8'h00;
            16'd26246: data <= 8'h1F;
            16'd26247: data <= 8'h00;
            16'd26248: data <= 8'h1F;
            16'd26249: data <= 8'h00;
            16'd26250: data <= 8'h1F;
            16'd26251: data <= 8'h00;
            16'd26252: data <= 8'h1F;
            16'd26253: data <= 8'h00;
            16'd26254: data <= 8'h1F;
            16'd26255: data <= 8'h00;
            16'd26256: data <= 8'h1F;
            16'd26257: data <= 8'h00;
            16'd26258: data <= 8'h1F;
            16'd26259: data <= 8'h00;
            16'd26260: data <= 8'h1F;
            16'd26261: data <= 8'h00;
            16'd26262: data <= 8'h1F;
            16'd26263: data <= 8'h00;
            16'd26264: data <= 8'h1F;
            16'd26265: data <= 8'h00;
            16'd26266: data <= 8'h1F;
            16'd26267: data <= 8'h00;
            16'd26268: data <= 8'h1F;
            16'd26269: data <= 8'h00;
            16'd26270: data <= 8'h1F;
            16'd26271: data <= 8'h00;
            16'd26272: data <= 8'h1F;
            16'd26273: data <= 8'h00;
            16'd26274: data <= 8'h1F;
            16'd26275: data <= 8'h00;
            16'd26276: data <= 8'h1F;
            16'd26277: data <= 8'h00;
            16'd26278: data <= 8'h1F;
            16'd26279: data <= 8'h00;
            16'd26280: data <= 8'hFF;
            16'd26281: data <= 8'hFF;
            16'd26282: data <= 8'h1F;
            16'd26283: data <= 8'h00;
            16'd26284: data <= 8'h1F;
            16'd26285: data <= 8'h00;
            16'd26286: data <= 8'h1F;
            16'd26287: data <= 8'h00;
            16'd26288: data <= 8'h1F;
            16'd26289: data <= 8'h00;
            16'd26290: data <= 8'h1F;
            16'd26291: data <= 8'h00;
            16'd26292: data <= 8'h1F;
            16'd26293: data <= 8'h00;
            16'd26294: data <= 8'h1F;
            16'd26295: data <= 8'h00;
            16'd26296: data <= 8'h1F;
            16'd26297: data <= 8'h00;
            16'd26298: data <= 8'h1F;
            16'd26299: data <= 8'h00;
            16'd26300: data <= 8'h1F;
            16'd26301: data <= 8'h00;
            16'd26302: data <= 8'h1F;
            16'd26303: data <= 8'h00;
            16'd26304: data <= 8'h1F;
            16'd26305: data <= 8'h00;
            16'd26306: data <= 8'h1F;
            16'd26307: data <= 8'h00;
            16'd26308: data <= 8'h1F;
            16'd26309: data <= 8'h00;
            16'd26310: data <= 8'h1F;
            16'd26311: data <= 8'h00;
            16'd26312: data <= 8'h1F;
            16'd26313: data <= 8'h00;
            16'd26314: data <= 8'h1F;
            16'd26315: data <= 8'h00;
            16'd26316: data <= 8'h1F;
            16'd26317: data <= 8'h00;
            16'd26318: data <= 8'h1F;
            16'd26319: data <= 8'h00;
            16'd26320: data <= 8'hFF;
            16'd26321: data <= 8'hFF;
            16'd26322: data <= 8'h1F;
            16'd26323: data <= 8'h00;
            16'd26324: data <= 8'h1F;
            16'd26325: data <= 8'h00;
            16'd26326: data <= 8'h1F;
            16'd26327: data <= 8'h00;
            16'd26328: data <= 8'h1F;
            16'd26329: data <= 8'h00;
            16'd26330: data <= 8'h1F;
            16'd26331: data <= 8'h00;
            16'd26332: data <= 8'h1F;
            16'd26333: data <= 8'h00;
            16'd26334: data <= 8'h1F;
            16'd26335: data <= 8'h00;
            16'd26336: data <= 8'h1F;
            16'd26337: data <= 8'h00;
            16'd26338: data <= 8'h1F;
            16'd26339: data <= 8'h00;
            16'd26340: data <= 8'h1F;
            16'd26341: data <= 8'h00;
            16'd26342: data <= 8'h1F;
            16'd26343: data <= 8'h00;
            16'd26344: data <= 8'h1F;
            16'd26345: data <= 8'h00;
            16'd26346: data <= 8'h1F;
            16'd26347: data <= 8'h00;
            16'd26348: data <= 8'h1F;
            16'd26349: data <= 8'h00;
            16'd26350: data <= 8'h1F;
            16'd26351: data <= 8'h00;
            16'd26352: data <= 8'h1F;
            16'd26353: data <= 8'h00;
            16'd26354: data <= 8'h1F;
            16'd26355: data <= 8'h00;
            16'd26356: data <= 8'h1F;
            16'd26357: data <= 8'h00;
            16'd26358: data <= 8'h1F;
            16'd26359: data <= 8'h00;
            16'd26360: data <= 8'hFF;
            16'd26361: data <= 8'hFF;
            16'd26362: data <= 8'h1F;
            16'd26363: data <= 8'h00;
            16'd26364: data <= 8'h1F;
            16'd26365: data <= 8'h00;
            16'd26366: data <= 8'h1F;
            16'd26367: data <= 8'h00;
            16'd26368: data <= 8'h1F;
            16'd26369: data <= 8'h00;
            16'd26370: data <= 8'h1F;
            16'd26371: data <= 8'h00;
            16'd26372: data <= 8'h1F;
            16'd26373: data <= 8'h00;
            16'd26374: data <= 8'h1F;
            16'd26375: data <= 8'h00;
            16'd26376: data <= 8'h1F;
            16'd26377: data <= 8'h00;
            16'd26378: data <= 8'h1F;
            16'd26379: data <= 8'h00;
            16'd26380: data <= 8'h1F;
            16'd26381: data <= 8'h00;
            16'd26382: data <= 8'h1F;
            16'd26383: data <= 8'h00;
            16'd26384: data <= 8'h1F;
            16'd26385: data <= 8'h00;
            16'd26386: data <= 8'h1F;
            16'd26387: data <= 8'h00;
            16'd26388: data <= 8'h1F;
            16'd26389: data <= 8'h00;
            16'd26390: data <= 8'h1F;
            16'd26391: data <= 8'h00;
            16'd26392: data <= 8'h1F;
            16'd26393: data <= 8'h00;
            16'd26394: data <= 8'h1F;
            16'd26395: data <= 8'h00;
            16'd26396: data <= 8'h1F;
            16'd26397: data <= 8'h00;
            16'd26398: data <= 8'h1F;
            16'd26399: data <= 8'h00;
            16'd26400: data <= 8'hFF;
            16'd26401: data <= 8'hFF;
            16'd26402: data <= 8'h1F;
            16'd26403: data <= 8'h00;
            16'd26404: data <= 8'h1F;
            16'd26405: data <= 8'h00;
            16'd26406: data <= 8'h1F;
            16'd26407: data <= 8'h00;
            16'd26408: data <= 8'h1F;
            16'd26409: data <= 8'h00;
            16'd26410: data <= 8'h1F;
            16'd26411: data <= 8'h00;
            16'd26412: data <= 8'h1F;
            16'd26413: data <= 8'h00;
            16'd26414: data <= 8'h1F;
            16'd26415: data <= 8'h00;
            16'd26416: data <= 8'h1F;
            16'd26417: data <= 8'h00;
            16'd26418: data <= 8'h1F;
            16'd26419: data <= 8'h00;
            16'd26420: data <= 8'h1F;
            16'd26421: data <= 8'h00;
            16'd26422: data <= 8'h1F;
            16'd26423: data <= 8'h00;
            16'd26424: data <= 8'h1F;
            16'd26425: data <= 8'h00;
            16'd26426: data <= 8'h1F;
            16'd26427: data <= 8'h00;
            16'd26428: data <= 8'h1F;
            16'd26429: data <= 8'h00;
            16'd26430: data <= 8'h1F;
            16'd26431: data <= 8'h00;
            16'd26432: data <= 8'h1F;
            16'd26433: data <= 8'h00;
            16'd26434: data <= 8'h1F;
            16'd26435: data <= 8'h00;
            16'd26436: data <= 8'h1F;
            16'd26437: data <= 8'h00;
            16'd26438: data <= 8'h1F;
            16'd26439: data <= 8'h00;
            16'd26440: data <= 8'hFF;
            16'd26441: data <= 8'hFF;
            16'd26442: data <= 8'h1F;
            16'd26443: data <= 8'h00;
            16'd26444: data <= 8'h1F;
            16'd26445: data <= 8'h00;
            16'd26446: data <= 8'h1F;
            16'd26447: data <= 8'h00;
            16'd26448: data <= 8'h1F;
            16'd26449: data <= 8'h00;
            16'd26450: data <= 8'h1F;
            16'd26451: data <= 8'h00;
            16'd26452: data <= 8'h1F;
            16'd26453: data <= 8'h00;
            16'd26454: data <= 8'h1F;
            16'd26455: data <= 8'h00;
            16'd26456: data <= 8'h1F;
            16'd26457: data <= 8'h00;
            16'd26458: data <= 8'h1F;
            16'd26459: data <= 8'h00;
            16'd26460: data <= 8'h1F;
            16'd26461: data <= 8'h00;
            16'd26462: data <= 8'h1F;
            16'd26463: data <= 8'h00;
            16'd26464: data <= 8'h1F;
            16'd26465: data <= 8'h00;
            16'd26466: data <= 8'h1F;
            16'd26467: data <= 8'h00;
            16'd26468: data <= 8'h1F;
            16'd26469: data <= 8'h00;
            16'd26470: data <= 8'h1F;
            16'd26471: data <= 8'h00;
            16'd26472: data <= 8'h1F;
            16'd26473: data <= 8'h00;
            16'd26474: data <= 8'h1F;
            16'd26475: data <= 8'h00;
            16'd26476: data <= 8'h1F;
            16'd26477: data <= 8'h00;
            16'd26478: data <= 8'h1F;
            16'd26479: data <= 8'h00;
            16'd26480: data <= 8'hFF;
            16'd26481: data <= 8'hFF;
            16'd26482: data <= 8'h1F;
            16'd26483: data <= 8'h00;
            16'd26484: data <= 8'h1F;
            16'd26485: data <= 8'h00;
            16'd26486: data <= 8'h1F;
            16'd26487: data <= 8'h00;
            16'd26488: data <= 8'h1F;
            16'd26489: data <= 8'h00;
            16'd26490: data <= 8'h1F;
            16'd26491: data <= 8'h00;
            16'd26492: data <= 8'h1F;
            16'd26493: data <= 8'h00;
            16'd26494: data <= 8'h1F;
            16'd26495: data <= 8'h00;
            16'd26496: data <= 8'h1F;
            16'd26497: data <= 8'h00;
            16'd26498: data <= 8'h1F;
            16'd26499: data <= 8'h00;
            16'd26500: data <= 8'h1F;
            16'd26501: data <= 8'h00;
            16'd26502: data <= 8'h1F;
            16'd26503: data <= 8'h00;
            16'd26504: data <= 8'h1F;
            16'd26505: data <= 8'h00;
            16'd26506: data <= 8'h1F;
            16'd26507: data <= 8'h00;
            16'd26508: data <= 8'h1F;
            16'd26509: data <= 8'h00;
            16'd26510: data <= 8'h1F;
            16'd26511: data <= 8'h00;
            16'd26512: data <= 8'h1F;
            16'd26513: data <= 8'h00;
            16'd26514: data <= 8'h1F;
            16'd26515: data <= 8'h00;
            16'd26516: data <= 8'h1F;
            16'd26517: data <= 8'h00;
            16'd26518: data <= 8'h1F;
            16'd26519: data <= 8'h00;
            16'd26520: data <= 8'hFF;
            16'd26521: data <= 8'hFF;
            16'd26522: data <= 8'h1F;
            16'd26523: data <= 8'h00;
            16'd26524: data <= 8'h1F;
            16'd26525: data <= 8'h00;
            16'd26526: data <= 8'h1F;
            16'd26527: data <= 8'h00;
            16'd26528: data <= 8'h1F;
            16'd26529: data <= 8'h00;
            16'd26530: data <= 8'h1F;
            16'd26531: data <= 8'h00;
            16'd26532: data <= 8'h1F;
            16'd26533: data <= 8'h00;
            16'd26534: data <= 8'h1F;
            16'd26535: data <= 8'h00;
            16'd26536: data <= 8'h1F;
            16'd26537: data <= 8'h00;
            16'd26538: data <= 8'h1F;
            16'd26539: data <= 8'h00;
            16'd26540: data <= 8'h1F;
            16'd26541: data <= 8'h00;
            16'd26542: data <= 8'h1F;
            16'd26543: data <= 8'h00;
            16'd26544: data <= 8'h1F;
            16'd26545: data <= 8'h00;
            16'd26546: data <= 8'h1F;
            16'd26547: data <= 8'h00;
            16'd26548: data <= 8'h1F;
            16'd26549: data <= 8'h00;
            16'd26550: data <= 8'h1F;
            16'd26551: data <= 8'h00;
            16'd26552: data <= 8'h1F;
            16'd26553: data <= 8'h00;
            16'd26554: data <= 8'h1F;
            16'd26555: data <= 8'h00;
            16'd26556: data <= 8'h1F;
            16'd26557: data <= 8'h00;
            16'd26558: data <= 8'h1F;
            16'd26559: data <= 8'h00;
            16'd26560: data <= 8'hFF;
            16'd26561: data <= 8'hFF;
            16'd26562: data <= 8'h1F;
            16'd26563: data <= 8'h00;
            16'd26564: data <= 8'h1F;
            16'd26565: data <= 8'h00;
            16'd26566: data <= 8'h1F;
            16'd26567: data <= 8'h00;
            16'd26568: data <= 8'h1F;
            16'd26569: data <= 8'h00;
            16'd26570: data <= 8'h1F;
            16'd26571: data <= 8'h00;
            16'd26572: data <= 8'h1F;
            16'd26573: data <= 8'h00;
            16'd26574: data <= 8'h1F;
            16'd26575: data <= 8'h00;
            16'd26576: data <= 8'h1F;
            16'd26577: data <= 8'h00;
            16'd26578: data <= 8'h1F;
            16'd26579: data <= 8'h00;
            16'd26580: data <= 8'h1F;
            16'd26581: data <= 8'h00;
            16'd26582: data <= 8'h1F;
            16'd26583: data <= 8'h00;
            16'd26584: data <= 8'h1F;
            16'd26585: data <= 8'h00;
            16'd26586: data <= 8'h1F;
            16'd26587: data <= 8'h00;
            16'd26588: data <= 8'h1F;
            16'd26589: data <= 8'h00;
            16'd26590: data <= 8'h1F;
            16'd26591: data <= 8'h00;
            16'd26592: data <= 8'h1F;
            16'd26593: data <= 8'h00;
            16'd26594: data <= 8'h1F;
            16'd26595: data <= 8'h00;
            16'd26596: data <= 8'h1F;
            16'd26597: data <= 8'h00;
            16'd26598: data <= 8'h1F;
            16'd26599: data <= 8'h00;
            16'd26600: data <= 8'hFF;
            16'd26601: data <= 8'hFF;
            16'd26602: data <= 8'h1F;
            16'd26603: data <= 8'h00;
            16'd26604: data <= 8'h1F;
            16'd26605: data <= 8'h00;
            16'd26606: data <= 8'h1F;
            16'd26607: data <= 8'h00;
            16'd26608: data <= 8'h1F;
            16'd26609: data <= 8'h00;
            16'd26610: data <= 8'h1F;
            16'd26611: data <= 8'h00;
            16'd26612: data <= 8'h1F;
            16'd26613: data <= 8'h00;
            16'd26614: data <= 8'h1F;
            16'd26615: data <= 8'h00;
            16'd26616: data <= 8'h1F;
            16'd26617: data <= 8'h00;
            16'd26618: data <= 8'h1F;
            16'd26619: data <= 8'h00;
            16'd26620: data <= 8'h1F;
            16'd26621: data <= 8'h00;
            16'd26622: data <= 8'h1F;
            16'd26623: data <= 8'h00;
            16'd26624: data <= 8'h1F;
            16'd26625: data <= 8'h00;
            16'd26626: data <= 8'h1F;
            16'd26627: data <= 8'h00;
            16'd26628: data <= 8'h1F;
            16'd26629: data <= 8'h00;
            16'd26630: data <= 8'h1F;
            16'd26631: data <= 8'h00;
            16'd26632: data <= 8'h1F;
            16'd26633: data <= 8'h00;
            16'd26634: data <= 8'h1F;
            16'd26635: data <= 8'h00;
            16'd26636: data <= 8'h1F;
            16'd26637: data <= 8'h00;
            16'd26638: data <= 8'h1F;
            16'd26639: data <= 8'h00;
            16'd26640: data <= 8'hFF;
            16'd26641: data <= 8'hFF;
            16'd26642: data <= 8'h1F;
            16'd26643: data <= 8'h00;
            16'd26644: data <= 8'h1F;
            16'd26645: data <= 8'h00;
            16'd26646: data <= 8'h1F;
            16'd26647: data <= 8'h00;
            16'd26648: data <= 8'h1F;
            16'd26649: data <= 8'h00;
            16'd26650: data <= 8'h1F;
            16'd26651: data <= 8'h00;
            16'd26652: data <= 8'h1F;
            16'd26653: data <= 8'h00;
            16'd26654: data <= 8'h1F;
            16'd26655: data <= 8'h00;
            16'd26656: data <= 8'h1F;
            16'd26657: data <= 8'h00;
            16'd26658: data <= 8'h1F;
            16'd26659: data <= 8'h00;
            16'd26660: data <= 8'h1F;
            16'd26661: data <= 8'h00;
            16'd26662: data <= 8'h1F;
            16'd26663: data <= 8'h00;
            16'd26664: data <= 8'h1F;
            16'd26665: data <= 8'h00;
            16'd26666: data <= 8'h1F;
            16'd26667: data <= 8'h00;
            16'd26668: data <= 8'h1F;
            16'd26669: data <= 8'h00;
            16'd26670: data <= 8'h1F;
            16'd26671: data <= 8'h00;
            16'd26672: data <= 8'h1F;
            16'd26673: data <= 8'h00;
            16'd26674: data <= 8'h1F;
            16'd26675: data <= 8'h00;
            16'd26676: data <= 8'h1F;
            16'd26677: data <= 8'h00;
            16'd26678: data <= 8'h1F;
            16'd26679: data <= 8'h00;
            16'd26680: data <= 8'hFF;
            16'd26681: data <= 8'hFF;
            16'd26682: data <= 8'h1F;
            16'd26683: data <= 8'h00;
            16'd26684: data <= 8'h1F;
            16'd26685: data <= 8'h00;
            16'd26686: data <= 8'h1F;
            16'd26687: data <= 8'h00;
            16'd26688: data <= 8'h1F;
            16'd26689: data <= 8'h00;
            16'd26690: data <= 8'h1F;
            16'd26691: data <= 8'h00;
            16'd26692: data <= 8'h1F;
            16'd26693: data <= 8'h00;
            16'd26694: data <= 8'h1F;
            16'd26695: data <= 8'h00;
            16'd26696: data <= 8'h1F;
            16'd26697: data <= 8'h00;
            16'd26698: data <= 8'h1F;
            16'd26699: data <= 8'h00;
            16'd26700: data <= 8'h1F;
            16'd26701: data <= 8'h00;
            16'd26702: data <= 8'h1F;
            16'd26703: data <= 8'h00;
            16'd26704: data <= 8'h1F;
            16'd26705: data <= 8'h00;
            16'd26706: data <= 8'h1F;
            16'd26707: data <= 8'h00;
            16'd26708: data <= 8'h1F;
            16'd26709: data <= 8'h00;
            16'd26710: data <= 8'h1F;
            16'd26711: data <= 8'h00;
            16'd26712: data <= 8'h1F;
            16'd26713: data <= 8'h00;
            16'd26714: data <= 8'h1F;
            16'd26715: data <= 8'h00;
            16'd26716: data <= 8'h1F;
            16'd26717: data <= 8'h00;
            16'd26718: data <= 8'h1F;
            16'd26719: data <= 8'h00;
            16'd26720: data <= 8'hFF;
            16'd26721: data <= 8'hFF;
            16'd26722: data <= 8'h1F;
            16'd26723: data <= 8'h00;
            16'd26724: data <= 8'h1F;
            16'd26725: data <= 8'h00;
            16'd26726: data <= 8'h1F;
            16'd26727: data <= 8'h00;
            16'd26728: data <= 8'h1F;
            16'd26729: data <= 8'h00;
            16'd26730: data <= 8'h1F;
            16'd26731: data <= 8'h00;
            16'd26732: data <= 8'h1F;
            16'd26733: data <= 8'h00;
            16'd26734: data <= 8'h1F;
            16'd26735: data <= 8'h00;
            16'd26736: data <= 8'h1F;
            16'd26737: data <= 8'h00;
            16'd26738: data <= 8'h1F;
            16'd26739: data <= 8'h00;
            16'd26740: data <= 8'h1F;
            16'd26741: data <= 8'h00;
            16'd26742: data <= 8'h1F;
            16'd26743: data <= 8'h00;
            16'd26744: data <= 8'h1F;
            16'd26745: data <= 8'h00;
            16'd26746: data <= 8'h1F;
            16'd26747: data <= 8'h00;
            16'd26748: data <= 8'h1F;
            16'd26749: data <= 8'h00;
            16'd26750: data <= 8'h1F;
            16'd26751: data <= 8'h00;
            16'd26752: data <= 8'h1F;
            16'd26753: data <= 8'h00;
            16'd26754: data <= 8'h1F;
            16'd26755: data <= 8'h00;
            16'd26756: data <= 8'h1F;
            16'd26757: data <= 8'h00;
            16'd26758: data <= 8'h1F;
            16'd26759: data <= 8'h00;
            16'd26760: data <= 8'hFF;
            16'd26761: data <= 8'hFF;
            16'd26762: data <= 8'h1F;
            16'd26763: data <= 8'h00;
            16'd26764: data <= 8'h1F;
            16'd26765: data <= 8'h00;
            16'd26766: data <= 8'h1F;
            16'd26767: data <= 8'h00;
            16'd26768: data <= 8'h1F;
            16'd26769: data <= 8'h00;
            16'd26770: data <= 8'h1F;
            16'd26771: data <= 8'h00;
            16'd26772: data <= 8'h1F;
            16'd26773: data <= 8'h00;
            16'd26774: data <= 8'h1F;
            16'd26775: data <= 8'h00;
            16'd26776: data <= 8'h1F;
            16'd26777: data <= 8'h00;
            16'd26778: data <= 8'h1F;
            16'd26779: data <= 8'h00;
            16'd26780: data <= 8'h1F;
            16'd26781: data <= 8'h00;
            16'd26782: data <= 8'h1F;
            16'd26783: data <= 8'h00;
            16'd26784: data <= 8'h1F;
            16'd26785: data <= 8'h00;
            16'd26786: data <= 8'h1F;
            16'd26787: data <= 8'h00;
            16'd26788: data <= 8'h1F;
            16'd26789: data <= 8'h00;
            16'd26790: data <= 8'h1F;
            16'd26791: data <= 8'h00;
            16'd26792: data <= 8'h1F;
            16'd26793: data <= 8'h00;
            16'd26794: data <= 8'h1F;
            16'd26795: data <= 8'h00;
            16'd26796: data <= 8'h1F;
            16'd26797: data <= 8'h00;
            16'd26798: data <= 8'h1F;
            16'd26799: data <= 8'h00;
            16'd26800: data <= 8'hFF;
            16'd26801: data <= 8'hFF;
            16'd26802: data <= 8'h1F;
            16'd26803: data <= 8'h00;
            16'd26804: data <= 8'h1F;
            16'd26805: data <= 8'h00;
            16'd26806: data <= 8'h1F;
            16'd26807: data <= 8'h00;
            16'd26808: data <= 8'h1F;
            16'd26809: data <= 8'h00;
            16'd26810: data <= 8'h1F;
            16'd26811: data <= 8'h00;
            16'd26812: data <= 8'h1F;
            16'd26813: data <= 8'h00;
            16'd26814: data <= 8'h1F;
            16'd26815: data <= 8'h00;
            16'd26816: data <= 8'h1F;
            16'd26817: data <= 8'h00;
            16'd26818: data <= 8'h1F;
            16'd26819: data <= 8'h00;
            16'd26820: data <= 8'h1F;
            16'd26821: data <= 8'h00;
            16'd26822: data <= 8'h1F;
            16'd26823: data <= 8'h00;
            16'd26824: data <= 8'h1F;
            16'd26825: data <= 8'h00;
            16'd26826: data <= 8'h1F;
            16'd26827: data <= 8'h00;
            16'd26828: data <= 8'h1F;
            16'd26829: data <= 8'h00;
            16'd26830: data <= 8'h1F;
            16'd26831: data <= 8'h00;
            16'd26832: data <= 8'h1F;
            16'd26833: data <= 8'h00;
            16'd26834: data <= 8'h1F;
            16'd26835: data <= 8'h00;
            16'd26836: data <= 8'h1F;
            16'd26837: data <= 8'h00;
            16'd26838: data <= 8'h1F;
            16'd26839: data <= 8'h00;
            16'd26840: data <= 8'hFF;
            16'd26841: data <= 8'hFF;
            16'd26842: data <= 8'h1F;
            16'd26843: data <= 8'h00;
            16'd26844: data <= 8'h1F;
            16'd26845: data <= 8'h00;
            16'd26846: data <= 8'h1F;
            16'd26847: data <= 8'h00;
            16'd26848: data <= 8'h1F;
            16'd26849: data <= 8'h00;
            16'd26850: data <= 8'h1F;
            16'd26851: data <= 8'h00;
            16'd26852: data <= 8'h1F;
            16'd26853: data <= 8'h00;
            16'd26854: data <= 8'h1F;
            16'd26855: data <= 8'h00;
            16'd26856: data <= 8'h1F;
            16'd26857: data <= 8'h00;
            16'd26858: data <= 8'h1F;
            16'd26859: data <= 8'h00;
            16'd26860: data <= 8'h1F;
            16'd26861: data <= 8'h00;
            16'd26862: data <= 8'h1F;
            16'd26863: data <= 8'h00;
            16'd26864: data <= 8'h1F;
            16'd26865: data <= 8'h00;
            16'd26866: data <= 8'h1F;
            16'd26867: data <= 8'h00;
            16'd26868: data <= 8'h1F;
            16'd26869: data <= 8'h00;
            16'd26870: data <= 8'h1F;
            16'd26871: data <= 8'h00;
            16'd26872: data <= 8'h1F;
            16'd26873: data <= 8'h00;
            16'd26874: data <= 8'h1F;
            16'd26875: data <= 8'h00;
            16'd26876: data <= 8'h1F;
            16'd26877: data <= 8'h00;
            16'd26878: data <= 8'h1F;
            16'd26879: data <= 8'h00;
            16'd26880: data <= 8'hFF;
            16'd26881: data <= 8'hFF;
            16'd26882: data <= 8'h1F;
            16'd26883: data <= 8'h00;
            16'd26884: data <= 8'h1F;
            16'd26885: data <= 8'h00;
            16'd26886: data <= 8'h1F;
            16'd26887: data <= 8'h00;
            16'd26888: data <= 8'h1F;
            16'd26889: data <= 8'h00;
            16'd26890: data <= 8'h1F;
            16'd26891: data <= 8'h00;
            16'd26892: data <= 8'h1F;
            16'd26893: data <= 8'h00;
            16'd26894: data <= 8'h1F;
            16'd26895: data <= 8'h00;
            16'd26896: data <= 8'h1F;
            16'd26897: data <= 8'h00;
            16'd26898: data <= 8'h1F;
            16'd26899: data <= 8'h00;
            16'd26900: data <= 8'h1F;
            16'd26901: data <= 8'h00;
            16'd26902: data <= 8'h1F;
            16'd26903: data <= 8'h00;
            16'd26904: data <= 8'h1F;
            16'd26905: data <= 8'h00;
            16'd26906: data <= 8'h1F;
            16'd26907: data <= 8'h00;
            16'd26908: data <= 8'h1F;
            16'd26909: data <= 8'h00;
            16'd26910: data <= 8'h1F;
            16'd26911: data <= 8'h00;
            16'd26912: data <= 8'h1F;
            16'd26913: data <= 8'h00;
            16'd26914: data <= 8'h1F;
            16'd26915: data <= 8'h00;
            16'd26916: data <= 8'h1F;
            16'd26917: data <= 8'h00;
            16'd26918: data <= 8'h1F;
            16'd26919: data <= 8'h00;
            16'd26920: data <= 8'hFF;
            16'd26921: data <= 8'hFF;
            16'd26922: data <= 8'h1F;
            16'd26923: data <= 8'h00;
            16'd26924: data <= 8'h1F;
            16'd26925: data <= 8'h00;
            16'd26926: data <= 8'h1F;
            16'd26927: data <= 8'h00;
            16'd26928: data <= 8'h1F;
            16'd26929: data <= 8'h00;
            16'd26930: data <= 8'h1F;
            16'd26931: data <= 8'h00;
            16'd26932: data <= 8'h1F;
            16'd26933: data <= 8'h00;
            16'd26934: data <= 8'h1F;
            16'd26935: data <= 8'h00;
            16'd26936: data <= 8'h1F;
            16'd26937: data <= 8'h00;
            16'd26938: data <= 8'h1F;
            16'd26939: data <= 8'h00;
            16'd26940: data <= 8'h1F;
            16'd26941: data <= 8'h00;
            16'd26942: data <= 8'h1F;
            16'd26943: data <= 8'h00;
            16'd26944: data <= 8'h1F;
            16'd26945: data <= 8'h00;
            16'd26946: data <= 8'h1F;
            16'd26947: data <= 8'h00;
            16'd26948: data <= 8'h1F;
            16'd26949: data <= 8'h00;
            16'd26950: data <= 8'h1F;
            16'd26951: data <= 8'h00;
            16'd26952: data <= 8'h1F;
            16'd26953: data <= 8'h00;
            16'd26954: data <= 8'h1F;
            16'd26955: data <= 8'h00;
            16'd26956: data <= 8'h1F;
            16'd26957: data <= 8'h00;
            16'd26958: data <= 8'h1F;
            16'd26959: data <= 8'h00;
            16'd26960: data <= 8'hFF;
            16'd26961: data <= 8'hFF;
            16'd26962: data <= 8'h1F;
            16'd26963: data <= 8'h00;
            16'd26964: data <= 8'h1F;
            16'd26965: data <= 8'h00;
            16'd26966: data <= 8'h1F;
            16'd26967: data <= 8'h00;
            16'd26968: data <= 8'h1F;
            16'd26969: data <= 8'h00;
            16'd26970: data <= 8'h1F;
            16'd26971: data <= 8'h00;
            16'd26972: data <= 8'h1F;
            16'd26973: data <= 8'h00;
            16'd26974: data <= 8'h1F;
            16'd26975: data <= 8'h00;
            16'd26976: data <= 8'h1F;
            16'd26977: data <= 8'h00;
            16'd26978: data <= 8'h1F;
            16'd26979: data <= 8'h00;
            16'd26980: data <= 8'h1F;
            16'd26981: data <= 8'h00;
            16'd26982: data <= 8'h1F;
            16'd26983: data <= 8'h00;
            16'd26984: data <= 8'h1F;
            16'd26985: data <= 8'h00;
            16'd26986: data <= 8'h1F;
            16'd26987: data <= 8'h00;
            16'd26988: data <= 8'h1F;
            16'd26989: data <= 8'h00;
            16'd26990: data <= 8'h1F;
            16'd26991: data <= 8'h00;
            16'd26992: data <= 8'h1F;
            16'd26993: data <= 8'h00;
            16'd26994: data <= 8'h1F;
            16'd26995: data <= 8'h00;
            16'd26996: data <= 8'h1F;
            16'd26997: data <= 8'h00;
            16'd26998: data <= 8'h1F;
            16'd26999: data <= 8'h00;
            16'd27000: data <= 8'hFF;
            16'd27001: data <= 8'hFF;
            16'd27002: data <= 8'h1F;
            16'd27003: data <= 8'h00;
            16'd27004: data <= 8'h1F;
            16'd27005: data <= 8'h00;
            16'd27006: data <= 8'h1F;
            16'd27007: data <= 8'h00;
            16'd27008: data <= 8'h1F;
            16'd27009: data <= 8'h00;
            16'd27010: data <= 8'h1F;
            16'd27011: data <= 8'h00;
            16'd27012: data <= 8'h1F;
            16'd27013: data <= 8'h00;
            16'd27014: data <= 8'h1F;
            16'd27015: data <= 8'h00;
            16'd27016: data <= 8'h1F;
            16'd27017: data <= 8'h00;
            16'd27018: data <= 8'h1F;
            16'd27019: data <= 8'h00;
            16'd27020: data <= 8'h1F;
            16'd27021: data <= 8'h00;
            16'd27022: data <= 8'h1F;
            16'd27023: data <= 8'h00;
            16'd27024: data <= 8'h1F;
            16'd27025: data <= 8'h00;
            16'd27026: data <= 8'h1F;
            16'd27027: data <= 8'h00;
            16'd27028: data <= 8'h1F;
            16'd27029: data <= 8'h00;
            16'd27030: data <= 8'h1F;
            16'd27031: data <= 8'h00;
            16'd27032: data <= 8'h1F;
            16'd27033: data <= 8'h00;
            16'd27034: data <= 8'h1F;
            16'd27035: data <= 8'h00;
            16'd27036: data <= 8'h1F;
            16'd27037: data <= 8'h00;
            16'd27038: data <= 8'h1F;
            16'd27039: data <= 8'h00;
            16'd27040: data <= 8'hFF;
            16'd27041: data <= 8'hFF;
            16'd27042: data <= 8'h1F;
            16'd27043: data <= 8'h00;
            16'd27044: data <= 8'h1F;
            16'd27045: data <= 8'h00;
            16'd27046: data <= 8'h1F;
            16'd27047: data <= 8'h00;
            16'd27048: data <= 8'h1F;
            16'd27049: data <= 8'h00;
            16'd27050: data <= 8'h1F;
            16'd27051: data <= 8'h00;
            16'd27052: data <= 8'h1F;
            16'd27053: data <= 8'h00;
            16'd27054: data <= 8'h1F;
            16'd27055: data <= 8'h00;
            16'd27056: data <= 8'h1F;
            16'd27057: data <= 8'h00;
            16'd27058: data <= 8'h1F;
            16'd27059: data <= 8'h00;
            16'd27060: data <= 8'h1F;
            16'd27061: data <= 8'h00;
            16'd27062: data <= 8'h1F;
            16'd27063: data <= 8'h00;
            16'd27064: data <= 8'h1F;
            16'd27065: data <= 8'h00;
            16'd27066: data <= 8'h1F;
            16'd27067: data <= 8'h00;
            16'd27068: data <= 8'h1F;
            16'd27069: data <= 8'h00;
            16'd27070: data <= 8'h1F;
            16'd27071: data <= 8'h00;
            16'd27072: data <= 8'h1F;
            16'd27073: data <= 8'h00;
            16'd27074: data <= 8'h1F;
            16'd27075: data <= 8'h00;
            16'd27076: data <= 8'h1F;
            16'd27077: data <= 8'h00;
            16'd27078: data <= 8'h1F;
            16'd27079: data <= 8'h00;
            16'd27080: data <= 8'hFF;
            16'd27081: data <= 8'hFF;
            16'd27082: data <= 8'h1F;
            16'd27083: data <= 8'h00;
            16'd27084: data <= 8'h1F;
            16'd27085: data <= 8'h00;
            16'd27086: data <= 8'h1F;
            16'd27087: data <= 8'h00;
            16'd27088: data <= 8'h1F;
            16'd27089: data <= 8'h00;
            16'd27090: data <= 8'h1F;
            16'd27091: data <= 8'h00;
            16'd27092: data <= 8'h1F;
            16'd27093: data <= 8'h00;
            16'd27094: data <= 8'h1F;
            16'd27095: data <= 8'h00;
            16'd27096: data <= 8'h1F;
            16'd27097: data <= 8'h00;
            16'd27098: data <= 8'h1F;
            16'd27099: data <= 8'h00;
            16'd27100: data <= 8'h1F;
            16'd27101: data <= 8'h00;
            16'd27102: data <= 8'h1F;
            16'd27103: data <= 8'h00;
            16'd27104: data <= 8'h1F;
            16'd27105: data <= 8'h00;
            16'd27106: data <= 8'h1F;
            16'd27107: data <= 8'h00;
            16'd27108: data <= 8'h1F;
            16'd27109: data <= 8'h00;
            16'd27110: data <= 8'h1F;
            16'd27111: data <= 8'h00;
            16'd27112: data <= 8'h1F;
            16'd27113: data <= 8'h00;
            16'd27114: data <= 8'h1F;
            16'd27115: data <= 8'h00;
            16'd27116: data <= 8'h1F;
            16'd27117: data <= 8'h00;
            16'd27118: data <= 8'h1F;
            16'd27119: data <= 8'h00;
            16'd27120: data <= 8'hFF;
            16'd27121: data <= 8'hFF;
            16'd27122: data <= 8'h1F;
            16'd27123: data <= 8'h00;
            16'd27124: data <= 8'h1F;
            16'd27125: data <= 8'h00;
            16'd27126: data <= 8'h1F;
            16'd27127: data <= 8'h00;
            16'd27128: data <= 8'h1F;
            16'd27129: data <= 8'h00;
            16'd27130: data <= 8'h1F;
            16'd27131: data <= 8'h00;
            16'd27132: data <= 8'h1F;
            16'd27133: data <= 8'h00;
            16'd27134: data <= 8'h1F;
            16'd27135: data <= 8'h00;
            16'd27136: data <= 8'h1F;
            16'd27137: data <= 8'h00;
            16'd27138: data <= 8'h1F;
            16'd27139: data <= 8'h00;
            16'd27140: data <= 8'h1F;
            16'd27141: data <= 8'h00;
            16'd27142: data <= 8'h1F;
            16'd27143: data <= 8'h00;
            16'd27144: data <= 8'h1F;
            16'd27145: data <= 8'h00;
            16'd27146: data <= 8'h1F;
            16'd27147: data <= 8'h00;
            16'd27148: data <= 8'h1F;
            16'd27149: data <= 8'h00;
            16'd27150: data <= 8'h1F;
            16'd27151: data <= 8'h00;
            16'd27152: data <= 8'h1F;
            16'd27153: data <= 8'h00;
            16'd27154: data <= 8'h1F;
            16'd27155: data <= 8'h00;
            16'd27156: data <= 8'h1F;
            16'd27157: data <= 8'h00;
            16'd27158: data <= 8'h1F;
            16'd27159: data <= 8'h00;
            16'd27160: data <= 8'hFF;
            16'd27161: data <= 8'hFF;
            16'd27162: data <= 8'h1F;
            16'd27163: data <= 8'h00;
            16'd27164: data <= 8'h1F;
            16'd27165: data <= 8'h00;
            16'd27166: data <= 8'h1F;
            16'd27167: data <= 8'h00;
            16'd27168: data <= 8'h1F;
            16'd27169: data <= 8'h00;
            16'd27170: data <= 8'h1F;
            16'd27171: data <= 8'h00;
            16'd27172: data <= 8'h1F;
            16'd27173: data <= 8'h00;
            16'd27174: data <= 8'h1F;
            16'd27175: data <= 8'h00;
            16'd27176: data <= 8'h1F;
            16'd27177: data <= 8'h00;
            16'd27178: data <= 8'h1F;
            16'd27179: data <= 8'h00;
            16'd27180: data <= 8'h1F;
            16'd27181: data <= 8'h00;
            16'd27182: data <= 8'h1F;
            16'd27183: data <= 8'h00;
            16'd27184: data <= 8'h1F;
            16'd27185: data <= 8'h00;
            16'd27186: data <= 8'h1F;
            16'd27187: data <= 8'h00;
            16'd27188: data <= 8'h1F;
            16'd27189: data <= 8'h00;
            16'd27190: data <= 8'h1F;
            16'd27191: data <= 8'h00;
            16'd27192: data <= 8'h1F;
            16'd27193: data <= 8'h00;
            16'd27194: data <= 8'h1F;
            16'd27195: data <= 8'h00;
            16'd27196: data <= 8'h1F;
            16'd27197: data <= 8'h00;
            16'd27198: data <= 8'h1F;
            16'd27199: data <= 8'h00;
            16'd27200: data <= 8'hFF;
            16'd27201: data <= 8'hFF;
            16'd27202: data <= 8'h1F;
            16'd27203: data <= 8'h00;
            16'd27204: data <= 8'h1F;
            16'd27205: data <= 8'h00;
            16'd27206: data <= 8'h1F;
            16'd27207: data <= 8'h00;
            16'd27208: data <= 8'h1F;
            16'd27209: data <= 8'h00;
            16'd27210: data <= 8'h1F;
            16'd27211: data <= 8'h00;
            16'd27212: data <= 8'h1F;
            16'd27213: data <= 8'h00;
            16'd27214: data <= 8'h1F;
            16'd27215: data <= 8'h00;
            16'd27216: data <= 8'h1F;
            16'd27217: data <= 8'h00;
            16'd27218: data <= 8'h1F;
            16'd27219: data <= 8'h00;
            16'd27220: data <= 8'h1F;
            16'd27221: data <= 8'h00;
            16'd27222: data <= 8'h1F;
            16'd27223: data <= 8'h00;
            16'd27224: data <= 8'h1F;
            16'd27225: data <= 8'h00;
            16'd27226: data <= 8'h1F;
            16'd27227: data <= 8'h00;
            16'd27228: data <= 8'h1F;
            16'd27229: data <= 8'h00;
            16'd27230: data <= 8'h1F;
            16'd27231: data <= 8'h00;
            16'd27232: data <= 8'h1F;
            16'd27233: data <= 8'h00;
            16'd27234: data <= 8'h1F;
            16'd27235: data <= 8'h00;
            16'd27236: data <= 8'h1F;
            16'd27237: data <= 8'h00;
            16'd27238: data <= 8'h1F;
            16'd27239: data <= 8'h00;
            16'd27240: data <= 8'hFF;
            16'd27241: data <= 8'hFF;
            16'd27242: data <= 8'h1F;
            16'd27243: data <= 8'h00;
            16'd27244: data <= 8'h1F;
            16'd27245: data <= 8'h00;
            16'd27246: data <= 8'h1F;
            16'd27247: data <= 8'h00;
            16'd27248: data <= 8'h1F;
            16'd27249: data <= 8'h00;
            16'd27250: data <= 8'h1F;
            16'd27251: data <= 8'h00;
            16'd27252: data <= 8'h1F;
            16'd27253: data <= 8'h00;
            16'd27254: data <= 8'h1F;
            16'd27255: data <= 8'h00;
            16'd27256: data <= 8'h1F;
            16'd27257: data <= 8'h00;
            16'd27258: data <= 8'h1F;
            16'd27259: data <= 8'h00;
            16'd27260: data <= 8'h1F;
            16'd27261: data <= 8'h00;
            16'd27262: data <= 8'h1F;
            16'd27263: data <= 8'h00;
            16'd27264: data <= 8'h1F;
            16'd27265: data <= 8'h00;
            16'd27266: data <= 8'h1F;
            16'd27267: data <= 8'h00;
            16'd27268: data <= 8'h1F;
            16'd27269: data <= 8'h00;
            16'd27270: data <= 8'h1F;
            16'd27271: data <= 8'h00;
            16'd27272: data <= 8'h1F;
            16'd27273: data <= 8'h00;
            16'd27274: data <= 8'h1F;
            16'd27275: data <= 8'h00;
            16'd27276: data <= 8'h1F;
            16'd27277: data <= 8'h00;
            16'd27278: data <= 8'h1F;
            16'd27279: data <= 8'h00;
            16'd27280: data <= 8'hFF;
            16'd27281: data <= 8'hFF;
            16'd27282: data <= 8'h1F;
            16'd27283: data <= 8'h00;
            16'd27284: data <= 8'h1F;
            16'd27285: data <= 8'h00;
            16'd27286: data <= 8'h1F;
            16'd27287: data <= 8'h00;
            16'd27288: data <= 8'h1F;
            16'd27289: data <= 8'h00;
            16'd27290: data <= 8'h1F;
            16'd27291: data <= 8'h00;
            16'd27292: data <= 8'h1F;
            16'd27293: data <= 8'h00;
            16'd27294: data <= 8'h1F;
            16'd27295: data <= 8'h00;
            16'd27296: data <= 8'h1F;
            16'd27297: data <= 8'h00;
            16'd27298: data <= 8'h1F;
            16'd27299: data <= 8'h00;
            16'd27300: data <= 8'h1F;
            16'd27301: data <= 8'h00;
            16'd27302: data <= 8'h1F;
            16'd27303: data <= 8'h00;
            16'd27304: data <= 8'h1F;
            16'd27305: data <= 8'h00;
            16'd27306: data <= 8'h1F;
            16'd27307: data <= 8'h00;
            16'd27308: data <= 8'h1F;
            16'd27309: data <= 8'h00;
            16'd27310: data <= 8'h1F;
            16'd27311: data <= 8'h00;
            16'd27312: data <= 8'h1F;
            16'd27313: data <= 8'h00;
            16'd27314: data <= 8'h1F;
            16'd27315: data <= 8'h00;
            16'd27316: data <= 8'h1F;
            16'd27317: data <= 8'h00;
            16'd27318: data <= 8'h1F;
            16'd27319: data <= 8'h00;
            16'd27320: data <= 8'hFF;
            16'd27321: data <= 8'hFF;
            16'd27322: data <= 8'h1F;
            16'd27323: data <= 8'h00;
            16'd27324: data <= 8'h1F;
            16'd27325: data <= 8'h00;
            16'd27326: data <= 8'h1F;
            16'd27327: data <= 8'h00;
            16'd27328: data <= 8'h1F;
            16'd27329: data <= 8'h00;
            16'd27330: data <= 8'h1F;
            16'd27331: data <= 8'h00;
            16'd27332: data <= 8'h1F;
            16'd27333: data <= 8'h00;
            16'd27334: data <= 8'h1F;
            16'd27335: data <= 8'h00;
            16'd27336: data <= 8'h1F;
            16'd27337: data <= 8'h00;
            16'd27338: data <= 8'h1F;
            16'd27339: data <= 8'h00;
            16'd27340: data <= 8'h1F;
            16'd27341: data <= 8'h00;
            16'd27342: data <= 8'h1F;
            16'd27343: data <= 8'h00;
            16'd27344: data <= 8'h1F;
            16'd27345: data <= 8'h00;
            16'd27346: data <= 8'h1F;
            16'd27347: data <= 8'h00;
            16'd27348: data <= 8'h1F;
            16'd27349: data <= 8'h00;
            16'd27350: data <= 8'h1F;
            16'd27351: data <= 8'h00;
            16'd27352: data <= 8'h1F;
            16'd27353: data <= 8'h00;
            16'd27354: data <= 8'h1F;
            16'd27355: data <= 8'h00;
            16'd27356: data <= 8'h1F;
            16'd27357: data <= 8'h00;
            16'd27358: data <= 8'h1F;
            16'd27359: data <= 8'h00;
            16'd27360: data <= 8'hFF;
            16'd27361: data <= 8'hFF;
            16'd27362: data <= 8'h1F;
            16'd27363: data <= 8'h00;
            16'd27364: data <= 8'h1F;
            16'd27365: data <= 8'h00;
            16'd27366: data <= 8'h1F;
            16'd27367: data <= 8'h00;
            16'd27368: data <= 8'h1F;
            16'd27369: data <= 8'h00;
            16'd27370: data <= 8'h1F;
            16'd27371: data <= 8'h00;
            16'd27372: data <= 8'h1F;
            16'd27373: data <= 8'h00;
            16'd27374: data <= 8'h1F;
            16'd27375: data <= 8'h00;
            16'd27376: data <= 8'h1F;
            16'd27377: data <= 8'h00;
            16'd27378: data <= 8'h1F;
            16'd27379: data <= 8'h00;
            16'd27380: data <= 8'h1F;
            16'd27381: data <= 8'h00;
            16'd27382: data <= 8'h1F;
            16'd27383: data <= 8'h00;
            16'd27384: data <= 8'h1F;
            16'd27385: data <= 8'h00;
            16'd27386: data <= 8'h1F;
            16'd27387: data <= 8'h00;
            16'd27388: data <= 8'h1F;
            16'd27389: data <= 8'h00;
            16'd27390: data <= 8'h1F;
            16'd27391: data <= 8'h00;
            16'd27392: data <= 8'h1F;
            16'd27393: data <= 8'h00;
            16'd27394: data <= 8'h1F;
            16'd27395: data <= 8'h00;
            16'd27396: data <= 8'h1F;
            16'd27397: data <= 8'h00;
            16'd27398: data <= 8'h1F;
            16'd27399: data <= 8'h00;
            16'd27400: data <= 8'hFF;
            16'd27401: data <= 8'hFF;
            16'd27402: data <= 8'h1F;
            16'd27403: data <= 8'h00;
            16'd27404: data <= 8'h1F;
            16'd27405: data <= 8'h00;
            16'd27406: data <= 8'h1F;
            16'd27407: data <= 8'h00;
            16'd27408: data <= 8'h1F;
            16'd27409: data <= 8'h00;
            16'd27410: data <= 8'h1F;
            16'd27411: data <= 8'h00;
            16'd27412: data <= 8'h1F;
            16'd27413: data <= 8'h00;
            16'd27414: data <= 8'h1F;
            16'd27415: data <= 8'h00;
            16'd27416: data <= 8'h1F;
            16'd27417: data <= 8'h00;
            16'd27418: data <= 8'h1F;
            16'd27419: data <= 8'h00;
            16'd27420: data <= 8'h1F;
            16'd27421: data <= 8'h00;
            16'd27422: data <= 8'h1F;
            16'd27423: data <= 8'h00;
            16'd27424: data <= 8'h1F;
            16'd27425: data <= 8'h00;
            16'd27426: data <= 8'h1F;
            16'd27427: data <= 8'h00;
            16'd27428: data <= 8'h1F;
            16'd27429: data <= 8'h00;
            16'd27430: data <= 8'h1F;
            16'd27431: data <= 8'h00;
            16'd27432: data <= 8'h1F;
            16'd27433: data <= 8'h00;
            16'd27434: data <= 8'h1F;
            16'd27435: data <= 8'h00;
            16'd27436: data <= 8'h1F;
            16'd27437: data <= 8'h00;
            16'd27438: data <= 8'h1F;
            16'd27439: data <= 8'h00;
            16'd27440: data <= 8'hFF;
            16'd27441: data <= 8'hFF;
            16'd27442: data <= 8'h1F;
            16'd27443: data <= 8'h00;
            16'd27444: data <= 8'h1F;
            16'd27445: data <= 8'h00;
            16'd27446: data <= 8'h1F;
            16'd27447: data <= 8'h00;
            16'd27448: data <= 8'h1F;
            16'd27449: data <= 8'h00;
            16'd27450: data <= 8'h1F;
            16'd27451: data <= 8'h00;
            16'd27452: data <= 8'h1F;
            16'd27453: data <= 8'h00;
            16'd27454: data <= 8'h1F;
            16'd27455: data <= 8'h00;
            16'd27456: data <= 8'h1F;
            16'd27457: data <= 8'h00;
            16'd27458: data <= 8'h1F;
            16'd27459: data <= 8'h00;
            16'd27460: data <= 8'h1F;
            16'd27461: data <= 8'h00;
            16'd27462: data <= 8'h1F;
            16'd27463: data <= 8'h00;
            16'd27464: data <= 8'h1F;
            16'd27465: data <= 8'h00;
            16'd27466: data <= 8'h1F;
            16'd27467: data <= 8'h00;
            16'd27468: data <= 8'h1F;
            16'd27469: data <= 8'h00;
            16'd27470: data <= 8'h1F;
            16'd27471: data <= 8'h00;
            16'd27472: data <= 8'h1F;
            16'd27473: data <= 8'h00;
            16'd27474: data <= 8'h1F;
            16'd27475: data <= 8'h00;
            16'd27476: data <= 8'h1F;
            16'd27477: data <= 8'h00;
            16'd27478: data <= 8'h1F;
            16'd27479: data <= 8'h00;
            16'd27480: data <= 8'hFF;
            16'd27481: data <= 8'hFF;
            16'd27482: data <= 8'h1F;
            16'd27483: data <= 8'h00;
            16'd27484: data <= 8'h1F;
            16'd27485: data <= 8'h00;
            16'd27486: data <= 8'h1F;
            16'd27487: data <= 8'h00;
            16'd27488: data <= 8'h1F;
            16'd27489: data <= 8'h00;
            16'd27490: data <= 8'h1F;
            16'd27491: data <= 8'h00;
            16'd27492: data <= 8'h1F;
            16'd27493: data <= 8'h00;
            16'd27494: data <= 8'h1F;
            16'd27495: data <= 8'h00;
            16'd27496: data <= 8'h1F;
            16'd27497: data <= 8'h00;
            16'd27498: data <= 8'h1F;
            16'd27499: data <= 8'h00;
            16'd27500: data <= 8'h1F;
            16'd27501: data <= 8'h00;
            16'd27502: data <= 8'h1F;
            16'd27503: data <= 8'h00;
            16'd27504: data <= 8'h1F;
            16'd27505: data <= 8'h00;
            16'd27506: data <= 8'h1F;
            16'd27507: data <= 8'h00;
            16'd27508: data <= 8'h1F;
            16'd27509: data <= 8'h00;
            16'd27510: data <= 8'h1F;
            16'd27511: data <= 8'h00;
            16'd27512: data <= 8'h1F;
            16'd27513: data <= 8'h00;
            16'd27514: data <= 8'h1F;
            16'd27515: data <= 8'h00;
            16'd27516: data <= 8'h1F;
            16'd27517: data <= 8'h00;
            16'd27518: data <= 8'h1F;
            16'd27519: data <= 8'h00;
            16'd27520: data <= 8'hFF;
            16'd27521: data <= 8'hFF;
            16'd27522: data <= 8'h1F;
            16'd27523: data <= 8'h00;
            16'd27524: data <= 8'h1F;
            16'd27525: data <= 8'h00;
            16'd27526: data <= 8'h1F;
            16'd27527: data <= 8'h00;
            16'd27528: data <= 8'h1F;
            16'd27529: data <= 8'h00;
            16'd27530: data <= 8'h1F;
            16'd27531: data <= 8'h00;
            16'd27532: data <= 8'h1F;
            16'd27533: data <= 8'h00;
            16'd27534: data <= 8'h1F;
            16'd27535: data <= 8'h00;
            16'd27536: data <= 8'h1F;
            16'd27537: data <= 8'h00;
            16'd27538: data <= 8'h1F;
            16'd27539: data <= 8'h00;
            16'd27540: data <= 8'h1F;
            16'd27541: data <= 8'h00;
            16'd27542: data <= 8'h1F;
            16'd27543: data <= 8'h00;
            16'd27544: data <= 8'h1F;
            16'd27545: data <= 8'h00;
            16'd27546: data <= 8'h1F;
            16'd27547: data <= 8'h00;
            16'd27548: data <= 8'h1F;
            16'd27549: data <= 8'h00;
            16'd27550: data <= 8'h1F;
            16'd27551: data <= 8'h00;
            16'd27552: data <= 8'h1F;
            16'd27553: data <= 8'h00;
            16'd27554: data <= 8'h1F;
            16'd27555: data <= 8'h00;
            16'd27556: data <= 8'h1F;
            16'd27557: data <= 8'h00;
            16'd27558: data <= 8'h1F;
            16'd27559: data <= 8'h00;
            16'd27560: data <= 8'hFF;
            16'd27561: data <= 8'hFF;
            16'd27562: data <= 8'h1F;
            16'd27563: data <= 8'h00;
            16'd27564: data <= 8'h1F;
            16'd27565: data <= 8'h00;
            16'd27566: data <= 8'h1F;
            16'd27567: data <= 8'h00;
            16'd27568: data <= 8'h1F;
            16'd27569: data <= 8'h00;
            16'd27570: data <= 8'h1F;
            16'd27571: data <= 8'h00;
            16'd27572: data <= 8'h1F;
            16'd27573: data <= 8'h00;
            16'd27574: data <= 8'h1F;
            16'd27575: data <= 8'h00;
            16'd27576: data <= 8'h1F;
            16'd27577: data <= 8'h00;
            16'd27578: data <= 8'h1F;
            16'd27579: data <= 8'h00;
            16'd27580: data <= 8'h1F;
            16'd27581: data <= 8'h00;
            16'd27582: data <= 8'h1F;
            16'd27583: data <= 8'h00;
            16'd27584: data <= 8'h1F;
            16'd27585: data <= 8'h00;
            16'd27586: data <= 8'h1F;
            16'd27587: data <= 8'h00;
            16'd27588: data <= 8'h1F;
            16'd27589: data <= 8'h00;
            16'd27590: data <= 8'h1F;
            16'd27591: data <= 8'h00;
            16'd27592: data <= 8'h1F;
            16'd27593: data <= 8'h00;
            16'd27594: data <= 8'h1F;
            16'd27595: data <= 8'h00;
            16'd27596: data <= 8'h1F;
            16'd27597: data <= 8'h00;
            16'd27598: data <= 8'h1F;
            16'd27599: data <= 8'h00;
            16'd27600: data <= 8'hFF;
            16'd27601: data <= 8'hFF;
            16'd27602: data <= 8'h1F;
            16'd27603: data <= 8'h00;
            16'd27604: data <= 8'h1F;
            16'd27605: data <= 8'h00;
            16'd27606: data <= 8'h1F;
            16'd27607: data <= 8'h00;
            16'd27608: data <= 8'h1F;
            16'd27609: data <= 8'h00;
            16'd27610: data <= 8'h1F;
            16'd27611: data <= 8'h00;
            16'd27612: data <= 8'h1F;
            16'd27613: data <= 8'h00;
            16'd27614: data <= 8'h1F;
            16'd27615: data <= 8'h00;
            16'd27616: data <= 8'h1F;
            16'd27617: data <= 8'h00;
            16'd27618: data <= 8'h1F;
            16'd27619: data <= 8'h00;
            16'd27620: data <= 8'h1F;
            16'd27621: data <= 8'h00;
            16'd27622: data <= 8'h1F;
            16'd27623: data <= 8'h00;
            16'd27624: data <= 8'h1F;
            16'd27625: data <= 8'h00;
            16'd27626: data <= 8'h1F;
            16'd27627: data <= 8'h00;
            16'd27628: data <= 8'h1F;
            16'd27629: data <= 8'h00;
            16'd27630: data <= 8'h1F;
            16'd27631: data <= 8'h00;
            16'd27632: data <= 8'h1F;
            16'd27633: data <= 8'h00;
            16'd27634: data <= 8'h1F;
            16'd27635: data <= 8'h00;
            16'd27636: data <= 8'h1F;
            16'd27637: data <= 8'h00;
            16'd27638: data <= 8'h1F;
            16'd27639: data <= 8'h00;
            16'd27640: data <= 8'hFF;
            16'd27641: data <= 8'hFF;
            16'd27642: data <= 8'h1F;
            16'd27643: data <= 8'h00;
            16'd27644: data <= 8'h1F;
            16'd27645: data <= 8'h00;
            16'd27646: data <= 8'h1F;
            16'd27647: data <= 8'h00;
            16'd27648: data <= 8'h1F;
            16'd27649: data <= 8'h00;
            16'd27650: data <= 8'h1F;
            16'd27651: data <= 8'h00;
            16'd27652: data <= 8'h1F;
            16'd27653: data <= 8'h00;
            16'd27654: data <= 8'h1F;
            16'd27655: data <= 8'h00;
            16'd27656: data <= 8'h1F;
            16'd27657: data <= 8'h00;
            16'd27658: data <= 8'h1F;
            16'd27659: data <= 8'h00;
            16'd27660: data <= 8'h1F;
            16'd27661: data <= 8'h00;
            16'd27662: data <= 8'h1F;
            16'd27663: data <= 8'h00;
            16'd27664: data <= 8'h1F;
            16'd27665: data <= 8'h00;
            16'd27666: data <= 8'h1F;
            16'd27667: data <= 8'h00;
            16'd27668: data <= 8'h1F;
            16'd27669: data <= 8'h00;
            16'd27670: data <= 8'h1F;
            16'd27671: data <= 8'h00;
            16'd27672: data <= 8'h1F;
            16'd27673: data <= 8'h00;
            16'd27674: data <= 8'h1F;
            16'd27675: data <= 8'h00;
            16'd27676: data <= 8'h1F;
            16'd27677: data <= 8'h00;
            16'd27678: data <= 8'h1F;
            16'd27679: data <= 8'h00;
            16'd27680: data <= 8'hFF;
            16'd27681: data <= 8'hFF;
            16'd27682: data <= 8'h1F;
            16'd27683: data <= 8'h00;
            16'd27684: data <= 8'h1F;
            16'd27685: data <= 8'h00;
            16'd27686: data <= 8'h1F;
            16'd27687: data <= 8'h00;
            16'd27688: data <= 8'h1F;
            16'd27689: data <= 8'h00;
            16'd27690: data <= 8'h1F;
            16'd27691: data <= 8'h00;
            16'd27692: data <= 8'h1F;
            16'd27693: data <= 8'h00;
            16'd27694: data <= 8'h1F;
            16'd27695: data <= 8'h00;
            16'd27696: data <= 8'h1F;
            16'd27697: data <= 8'h00;
            16'd27698: data <= 8'h1F;
            16'd27699: data <= 8'h00;
            16'd27700: data <= 8'h1F;
            16'd27701: data <= 8'h00;
            16'd27702: data <= 8'h1F;
            16'd27703: data <= 8'h00;
            16'd27704: data <= 8'h1F;
            16'd27705: data <= 8'h00;
            16'd27706: data <= 8'h1F;
            16'd27707: data <= 8'h00;
            16'd27708: data <= 8'h1F;
            16'd27709: data <= 8'h00;
            16'd27710: data <= 8'h1F;
            16'd27711: data <= 8'h00;
            16'd27712: data <= 8'h1F;
            16'd27713: data <= 8'h00;
            16'd27714: data <= 8'h1F;
            16'd27715: data <= 8'h00;
            16'd27716: data <= 8'h1F;
            16'd27717: data <= 8'h00;
            16'd27718: data <= 8'h1F;
            16'd27719: data <= 8'h00;
            16'd27720: data <= 8'hFF;
            16'd27721: data <= 8'hFF;
            16'd27722: data <= 8'h1F;
            16'd27723: data <= 8'h00;
            16'd27724: data <= 8'h1F;
            16'd27725: data <= 8'h00;
            16'd27726: data <= 8'h1F;
            16'd27727: data <= 8'h00;
            16'd27728: data <= 8'h1F;
            16'd27729: data <= 8'h00;
            16'd27730: data <= 8'h1F;
            16'd27731: data <= 8'h00;
            16'd27732: data <= 8'h1F;
            16'd27733: data <= 8'h00;
            16'd27734: data <= 8'h1F;
            16'd27735: data <= 8'h00;
            16'd27736: data <= 8'h1F;
            16'd27737: data <= 8'h00;
            16'd27738: data <= 8'h1F;
            16'd27739: data <= 8'h00;
            16'd27740: data <= 8'h1F;
            16'd27741: data <= 8'h00;
            16'd27742: data <= 8'h1F;
            16'd27743: data <= 8'h00;
            16'd27744: data <= 8'h1F;
            16'd27745: data <= 8'h00;
            16'd27746: data <= 8'h1F;
            16'd27747: data <= 8'h00;
            16'd27748: data <= 8'h1F;
            16'd27749: data <= 8'h00;
            16'd27750: data <= 8'h1F;
            16'd27751: data <= 8'h00;
            16'd27752: data <= 8'h1F;
            16'd27753: data <= 8'h00;
            16'd27754: data <= 8'h1F;
            16'd27755: data <= 8'h00;
            16'd27756: data <= 8'h1F;
            16'd27757: data <= 8'h00;
            16'd27758: data <= 8'h1F;
            16'd27759: data <= 8'h00;
            16'd27760: data <= 8'hFF;
            16'd27761: data <= 8'hFF;
            16'd27762: data <= 8'h1F;
            16'd27763: data <= 8'h00;
            16'd27764: data <= 8'h1F;
            16'd27765: data <= 8'h00;
            16'd27766: data <= 8'h1F;
            16'd27767: data <= 8'h00;
            16'd27768: data <= 8'h1F;
            16'd27769: data <= 8'h00;
            16'd27770: data <= 8'h1F;
            16'd27771: data <= 8'h00;
            16'd27772: data <= 8'h1F;
            16'd27773: data <= 8'h00;
            16'd27774: data <= 8'h1F;
            16'd27775: data <= 8'h00;
            16'd27776: data <= 8'h1F;
            16'd27777: data <= 8'h00;
            16'd27778: data <= 8'h1F;
            16'd27779: data <= 8'h00;
            16'd27780: data <= 8'h1F;
            16'd27781: data <= 8'h00;
            16'd27782: data <= 8'h1F;
            16'd27783: data <= 8'h00;
            16'd27784: data <= 8'h1F;
            16'd27785: data <= 8'h00;
            16'd27786: data <= 8'h1F;
            16'd27787: data <= 8'h00;
            16'd27788: data <= 8'h1F;
            16'd27789: data <= 8'h00;
            16'd27790: data <= 8'h1F;
            16'd27791: data <= 8'h00;
            16'd27792: data <= 8'h1F;
            16'd27793: data <= 8'h00;
            16'd27794: data <= 8'h1F;
            16'd27795: data <= 8'h00;
            16'd27796: data <= 8'h1F;
            16'd27797: data <= 8'h00;
            16'd27798: data <= 8'h1F;
            16'd27799: data <= 8'h00;
            16'd27800: data <= 8'hFF;
            16'd27801: data <= 8'hFF;
            16'd27802: data <= 8'h1F;
            16'd27803: data <= 8'h00;
            16'd27804: data <= 8'h1F;
            16'd27805: data <= 8'h00;
            16'd27806: data <= 8'h1F;
            16'd27807: data <= 8'h00;
            16'd27808: data <= 8'h1F;
            16'd27809: data <= 8'h00;
            16'd27810: data <= 8'h1F;
            16'd27811: data <= 8'h00;
            16'd27812: data <= 8'h1F;
            16'd27813: data <= 8'h00;
            16'd27814: data <= 8'h1F;
            16'd27815: data <= 8'h00;
            16'd27816: data <= 8'h1F;
            16'd27817: data <= 8'h00;
            16'd27818: data <= 8'h1F;
            16'd27819: data <= 8'h00;
            16'd27820: data <= 8'h1F;
            16'd27821: data <= 8'h00;
            16'd27822: data <= 8'h1F;
            16'd27823: data <= 8'h00;
            16'd27824: data <= 8'h1F;
            16'd27825: data <= 8'h00;
            16'd27826: data <= 8'h1F;
            16'd27827: data <= 8'h00;
            16'd27828: data <= 8'h1F;
            16'd27829: data <= 8'h00;
            16'd27830: data <= 8'h1F;
            16'd27831: data <= 8'h00;
            16'd27832: data <= 8'h1F;
            16'd27833: data <= 8'h00;
            16'd27834: data <= 8'h1F;
            16'd27835: data <= 8'h00;
            16'd27836: data <= 8'h1F;
            16'd27837: data <= 8'h00;
            16'd27838: data <= 8'h1F;
            16'd27839: data <= 8'h00;
            16'd27840: data <= 8'hFF;
            16'd27841: data <= 8'hFF;
            16'd27842: data <= 8'h1F;
            16'd27843: data <= 8'h00;
            16'd27844: data <= 8'h1F;
            16'd27845: data <= 8'h00;
            16'd27846: data <= 8'h1F;
            16'd27847: data <= 8'h00;
            16'd27848: data <= 8'h1F;
            16'd27849: data <= 8'h00;
            16'd27850: data <= 8'h1F;
            16'd27851: data <= 8'h00;
            16'd27852: data <= 8'h1F;
            16'd27853: data <= 8'h00;
            16'd27854: data <= 8'h1F;
            16'd27855: data <= 8'h00;
            16'd27856: data <= 8'h1F;
            16'd27857: data <= 8'h00;
            16'd27858: data <= 8'h1F;
            16'd27859: data <= 8'h00;
            16'd27860: data <= 8'h1F;
            16'd27861: data <= 8'h00;
            16'd27862: data <= 8'h1F;
            16'd27863: data <= 8'h00;
            16'd27864: data <= 8'h1F;
            16'd27865: data <= 8'h00;
            16'd27866: data <= 8'h1F;
            16'd27867: data <= 8'h00;
            16'd27868: data <= 8'h1F;
            16'd27869: data <= 8'h00;
            16'd27870: data <= 8'h1F;
            16'd27871: data <= 8'h00;
            16'd27872: data <= 8'h1F;
            16'd27873: data <= 8'h00;
            16'd27874: data <= 8'h1F;
            16'd27875: data <= 8'h00;
            16'd27876: data <= 8'h1F;
            16'd27877: data <= 8'h00;
            16'd27878: data <= 8'h1F;
            16'd27879: data <= 8'h00;
            16'd27880: data <= 8'hFF;
            16'd27881: data <= 8'hFF;
            16'd27882: data <= 8'h1F;
            16'd27883: data <= 8'h00;
            16'd27884: data <= 8'h1F;
            16'd27885: data <= 8'h00;
            16'd27886: data <= 8'h1F;
            16'd27887: data <= 8'h00;
            16'd27888: data <= 8'h1F;
            16'd27889: data <= 8'h00;
            16'd27890: data <= 8'h1F;
            16'd27891: data <= 8'h00;
            16'd27892: data <= 8'h1F;
            16'd27893: data <= 8'h00;
            16'd27894: data <= 8'h1F;
            16'd27895: data <= 8'h00;
            16'd27896: data <= 8'h1F;
            16'd27897: data <= 8'h00;
            16'd27898: data <= 8'h1F;
            16'd27899: data <= 8'h00;
            16'd27900: data <= 8'h1F;
            16'd27901: data <= 8'h00;
            16'd27902: data <= 8'h1F;
            16'd27903: data <= 8'h00;
            16'd27904: data <= 8'h1F;
            16'd27905: data <= 8'h00;
            16'd27906: data <= 8'h1F;
            16'd27907: data <= 8'h00;
            16'd27908: data <= 8'h1F;
            16'd27909: data <= 8'h00;
            16'd27910: data <= 8'h1F;
            16'd27911: data <= 8'h00;
            16'd27912: data <= 8'h1F;
            16'd27913: data <= 8'h00;
            16'd27914: data <= 8'h1F;
            16'd27915: data <= 8'h00;
            16'd27916: data <= 8'h1F;
            16'd27917: data <= 8'h00;
            16'd27918: data <= 8'h1F;
            16'd27919: data <= 8'h00;
            16'd27920: data <= 8'hFF;
            16'd27921: data <= 8'hFF;
            16'd27922: data <= 8'h1F;
            16'd27923: data <= 8'h00;
            16'd27924: data <= 8'h1F;
            16'd27925: data <= 8'h00;
            16'd27926: data <= 8'h1F;
            16'd27927: data <= 8'h00;
            16'd27928: data <= 8'h1F;
            16'd27929: data <= 8'h00;
            16'd27930: data <= 8'h1F;
            16'd27931: data <= 8'h00;
            16'd27932: data <= 8'h1F;
            16'd27933: data <= 8'h00;
            16'd27934: data <= 8'h1F;
            16'd27935: data <= 8'h00;
            16'd27936: data <= 8'h1F;
            16'd27937: data <= 8'h00;
            16'd27938: data <= 8'h1F;
            16'd27939: data <= 8'h00;
            16'd27940: data <= 8'h1F;
            16'd27941: data <= 8'h00;
            16'd27942: data <= 8'h1F;
            16'd27943: data <= 8'h00;
            16'd27944: data <= 8'h1F;
            16'd27945: data <= 8'h00;
            16'd27946: data <= 8'h1F;
            16'd27947: data <= 8'h00;
            16'd27948: data <= 8'h1F;
            16'd27949: data <= 8'h00;
            16'd27950: data <= 8'h1F;
            16'd27951: data <= 8'h00;
            16'd27952: data <= 8'h1F;
            16'd27953: data <= 8'h00;
            16'd27954: data <= 8'h1F;
            16'd27955: data <= 8'h00;
            16'd27956: data <= 8'h1F;
            16'd27957: data <= 8'h00;
            16'd27958: data <= 8'h1F;
            16'd27959: data <= 8'h00;
            16'd27960: data <= 8'hFF;
            16'd27961: data <= 8'hFF;
            16'd27962: data <= 8'h1F;
            16'd27963: data <= 8'h00;
            16'd27964: data <= 8'h1F;
            16'd27965: data <= 8'h00;
            16'd27966: data <= 8'h1F;
            16'd27967: data <= 8'h00;
            16'd27968: data <= 8'h1F;
            16'd27969: data <= 8'h00;
            16'd27970: data <= 8'h1F;
            16'd27971: data <= 8'h00;
            16'd27972: data <= 8'h1F;
            16'd27973: data <= 8'h00;
            16'd27974: data <= 8'h1F;
            16'd27975: data <= 8'h00;
            16'd27976: data <= 8'h1F;
            16'd27977: data <= 8'h00;
            16'd27978: data <= 8'h1F;
            16'd27979: data <= 8'h00;
            16'd27980: data <= 8'h1F;
            16'd27981: data <= 8'h00;
            16'd27982: data <= 8'h1F;
            16'd27983: data <= 8'h00;
            16'd27984: data <= 8'h1F;
            16'd27985: data <= 8'h00;
            16'd27986: data <= 8'h1F;
            16'd27987: data <= 8'h00;
            16'd27988: data <= 8'h1F;
            16'd27989: data <= 8'h00;
            16'd27990: data <= 8'h1F;
            16'd27991: data <= 8'h00;
            16'd27992: data <= 8'h1F;
            16'd27993: data <= 8'h00;
            16'd27994: data <= 8'h1F;
            16'd27995: data <= 8'h00;
            16'd27996: data <= 8'h1F;
            16'd27997: data <= 8'h00;
            16'd27998: data <= 8'h1F;
            16'd27999: data <= 8'h00;
            16'd28000: data <= 8'hFF;
            16'd28001: data <= 8'hFF;
            16'd28002: data <= 8'h1F;
            16'd28003: data <= 8'h00;
            16'd28004: data <= 8'h1F;
            16'd28005: data <= 8'h00;
            16'd28006: data <= 8'h1F;
            16'd28007: data <= 8'h00;
            16'd28008: data <= 8'h1F;
            16'd28009: data <= 8'h00;
            16'd28010: data <= 8'h1F;
            16'd28011: data <= 8'h00;
            16'd28012: data <= 8'h1F;
            16'd28013: data <= 8'h00;
            16'd28014: data <= 8'h1F;
            16'd28015: data <= 8'h00;
            16'd28016: data <= 8'h1F;
            16'd28017: data <= 8'h00;
            16'd28018: data <= 8'h1F;
            16'd28019: data <= 8'h00;
            16'd28020: data <= 8'h1F;
            16'd28021: data <= 8'h00;
            16'd28022: data <= 8'h1F;
            16'd28023: data <= 8'h00;
            16'd28024: data <= 8'h1F;
            16'd28025: data <= 8'h00;
            16'd28026: data <= 8'h1F;
            16'd28027: data <= 8'h00;
            16'd28028: data <= 8'h1F;
            16'd28029: data <= 8'h00;
            16'd28030: data <= 8'h1F;
            16'd28031: data <= 8'h00;
            16'd28032: data <= 8'h1F;
            16'd28033: data <= 8'h00;
            16'd28034: data <= 8'h1F;
            16'd28035: data <= 8'h00;
            16'd28036: data <= 8'h1F;
            16'd28037: data <= 8'h00;
            16'd28038: data <= 8'h1F;
            16'd28039: data <= 8'h00;
            16'd28040: data <= 8'hFF;
            16'd28041: data <= 8'hFF;
            16'd28042: data <= 8'h1F;
            16'd28043: data <= 8'h00;
            16'd28044: data <= 8'h1F;
            16'd28045: data <= 8'h00;
            16'd28046: data <= 8'h1F;
            16'd28047: data <= 8'h00;
            16'd28048: data <= 8'h1F;
            16'd28049: data <= 8'h00;
            16'd28050: data <= 8'h1F;
            16'd28051: data <= 8'h00;
            16'd28052: data <= 8'h1F;
            16'd28053: data <= 8'h00;
            16'd28054: data <= 8'h1F;
            16'd28055: data <= 8'h00;
            16'd28056: data <= 8'h1F;
            16'd28057: data <= 8'h00;
            16'd28058: data <= 8'h1F;
            16'd28059: data <= 8'h00;
            16'd28060: data <= 8'h1F;
            16'd28061: data <= 8'h00;
            16'd28062: data <= 8'h1F;
            16'd28063: data <= 8'h00;
            16'd28064: data <= 8'h1F;
            16'd28065: data <= 8'h00;
            16'd28066: data <= 8'h1F;
            16'd28067: data <= 8'h00;
            16'd28068: data <= 8'h1F;
            16'd28069: data <= 8'h00;
            16'd28070: data <= 8'h1F;
            16'd28071: data <= 8'h00;
            16'd28072: data <= 8'h1F;
            16'd28073: data <= 8'h00;
            16'd28074: data <= 8'h1F;
            16'd28075: data <= 8'h00;
            16'd28076: data <= 8'h1F;
            16'd28077: data <= 8'h00;
            16'd28078: data <= 8'h1F;
            16'd28079: data <= 8'h00;
            16'd28080: data <= 8'hFF;
            16'd28081: data <= 8'hFF;
            16'd28082: data <= 8'h1F;
            16'd28083: data <= 8'h00;
            16'd28084: data <= 8'h1F;
            16'd28085: data <= 8'h00;
            16'd28086: data <= 8'h1F;
            16'd28087: data <= 8'h00;
            16'd28088: data <= 8'h1F;
            16'd28089: data <= 8'h00;
            16'd28090: data <= 8'h1F;
            16'd28091: data <= 8'h00;
            16'd28092: data <= 8'h1F;
            16'd28093: data <= 8'h00;
            16'd28094: data <= 8'h1F;
            16'd28095: data <= 8'h00;
            16'd28096: data <= 8'h1F;
            16'd28097: data <= 8'h00;
            16'd28098: data <= 8'h1F;
            16'd28099: data <= 8'h00;
            16'd28100: data <= 8'h1F;
            16'd28101: data <= 8'h00;
            16'd28102: data <= 8'h1F;
            16'd28103: data <= 8'h00;
            16'd28104: data <= 8'h1F;
            16'd28105: data <= 8'h00;
            16'd28106: data <= 8'h1F;
            16'd28107: data <= 8'h00;
            16'd28108: data <= 8'h1F;
            16'd28109: data <= 8'h00;
            16'd28110: data <= 8'h1F;
            16'd28111: data <= 8'h00;
            16'd28112: data <= 8'h1F;
            16'd28113: data <= 8'h00;
            16'd28114: data <= 8'h1F;
            16'd28115: data <= 8'h00;
            16'd28116: data <= 8'h1F;
            16'd28117: data <= 8'h00;
            16'd28118: data <= 8'h1F;
            16'd28119: data <= 8'h00;
            16'd28120: data <= 8'hFF;
            16'd28121: data <= 8'hFF;
            16'd28122: data <= 8'h1F;
            16'd28123: data <= 8'h00;
            16'd28124: data <= 8'h1F;
            16'd28125: data <= 8'h00;
            16'd28126: data <= 8'h1F;
            16'd28127: data <= 8'h00;
            16'd28128: data <= 8'h1F;
            16'd28129: data <= 8'h00;
            16'd28130: data <= 8'h1F;
            16'd28131: data <= 8'h00;
            16'd28132: data <= 8'h1F;
            16'd28133: data <= 8'h00;
            16'd28134: data <= 8'h1F;
            16'd28135: data <= 8'h00;
            16'd28136: data <= 8'h1F;
            16'd28137: data <= 8'h00;
            16'd28138: data <= 8'h1F;
            16'd28139: data <= 8'h00;
            16'd28140: data <= 8'h1F;
            16'd28141: data <= 8'h00;
            16'd28142: data <= 8'h1F;
            16'd28143: data <= 8'h00;
            16'd28144: data <= 8'h1F;
            16'd28145: data <= 8'h00;
            16'd28146: data <= 8'h1F;
            16'd28147: data <= 8'h00;
            16'd28148: data <= 8'h1F;
            16'd28149: data <= 8'h00;
            16'd28150: data <= 8'h1F;
            16'd28151: data <= 8'h00;
            16'd28152: data <= 8'h1F;
            16'd28153: data <= 8'h00;
            16'd28154: data <= 8'h1F;
            16'd28155: data <= 8'h00;
            16'd28156: data <= 8'h1F;
            16'd28157: data <= 8'h00;
            16'd28158: data <= 8'h1F;
            16'd28159: data <= 8'h00;
            16'd28160: data <= 8'hFF;
            16'd28161: data <= 8'hFF;
            16'd28162: data <= 8'h1F;
            16'd28163: data <= 8'h00;
            16'd28164: data <= 8'h1F;
            16'd28165: data <= 8'h00;
            16'd28166: data <= 8'h1F;
            16'd28167: data <= 8'h00;
            16'd28168: data <= 8'h1F;
            16'd28169: data <= 8'h00;
            16'd28170: data <= 8'h1F;
            16'd28171: data <= 8'h00;
            16'd28172: data <= 8'h1F;
            16'd28173: data <= 8'h00;
            16'd28174: data <= 8'h1F;
            16'd28175: data <= 8'h00;
            16'd28176: data <= 8'h1F;
            16'd28177: data <= 8'h00;
            16'd28178: data <= 8'h1F;
            16'd28179: data <= 8'h00;
            16'd28180: data <= 8'h1F;
            16'd28181: data <= 8'h00;
            16'd28182: data <= 8'h1F;
            16'd28183: data <= 8'h00;
            16'd28184: data <= 8'h1F;
            16'd28185: data <= 8'h00;
            16'd28186: data <= 8'h1F;
            16'd28187: data <= 8'h00;
            16'd28188: data <= 8'h1F;
            16'd28189: data <= 8'h00;
            16'd28190: data <= 8'h1F;
            16'd28191: data <= 8'h00;
            16'd28192: data <= 8'h1F;
            16'd28193: data <= 8'h00;
            16'd28194: data <= 8'h1F;
            16'd28195: data <= 8'h00;
            16'd28196: data <= 8'h1F;
            16'd28197: data <= 8'h00;
            16'd28198: data <= 8'h1F;
            16'd28199: data <= 8'h00;
            16'd28200: data <= 8'hFF;
            16'd28201: data <= 8'hFF;
            16'd28202: data <= 8'h1F;
            16'd28203: data <= 8'h00;
            16'd28204: data <= 8'h1F;
            16'd28205: data <= 8'h00;
            16'd28206: data <= 8'h1F;
            16'd28207: data <= 8'h00;
            16'd28208: data <= 8'h1F;
            16'd28209: data <= 8'h00;
            16'd28210: data <= 8'h1F;
            16'd28211: data <= 8'h00;
            16'd28212: data <= 8'h1F;
            16'd28213: data <= 8'h00;
            16'd28214: data <= 8'h1F;
            16'd28215: data <= 8'h00;
            16'd28216: data <= 8'h1F;
            16'd28217: data <= 8'h00;
            16'd28218: data <= 8'h1F;
            16'd28219: data <= 8'h00;
            16'd28220: data <= 8'h1F;
            16'd28221: data <= 8'h00;
            16'd28222: data <= 8'h1F;
            16'd28223: data <= 8'h00;
            16'd28224: data <= 8'h1F;
            16'd28225: data <= 8'h00;
            16'd28226: data <= 8'h1F;
            16'd28227: data <= 8'h00;
            16'd28228: data <= 8'h1F;
            16'd28229: data <= 8'h00;
            16'd28230: data <= 8'h1F;
            16'd28231: data <= 8'h00;
            16'd28232: data <= 8'h1F;
            16'd28233: data <= 8'h00;
            16'd28234: data <= 8'h1F;
            16'd28235: data <= 8'h00;
            16'd28236: data <= 8'h1F;
            16'd28237: data <= 8'h00;
            16'd28238: data <= 8'h1F;
            16'd28239: data <= 8'h00;
            16'd28240: data <= 8'hFF;
            16'd28241: data <= 8'hFF;
            16'd28242: data <= 8'h1F;
            16'd28243: data <= 8'h00;
            16'd28244: data <= 8'h1F;
            16'd28245: data <= 8'h00;
            16'd28246: data <= 8'h1F;
            16'd28247: data <= 8'h00;
            16'd28248: data <= 8'h1F;
            16'd28249: data <= 8'h00;
            16'd28250: data <= 8'h1F;
            16'd28251: data <= 8'h00;
            16'd28252: data <= 8'h1F;
            16'd28253: data <= 8'h00;
            16'd28254: data <= 8'h1F;
            16'd28255: data <= 8'h00;
            16'd28256: data <= 8'h1F;
            16'd28257: data <= 8'h00;
            16'd28258: data <= 8'h1F;
            16'd28259: data <= 8'h00;
            16'd28260: data <= 8'h1F;
            16'd28261: data <= 8'h00;
            16'd28262: data <= 8'h1F;
            16'd28263: data <= 8'h00;
            16'd28264: data <= 8'h1F;
            16'd28265: data <= 8'h00;
            16'd28266: data <= 8'h1F;
            16'd28267: data <= 8'h00;
            16'd28268: data <= 8'h1F;
            16'd28269: data <= 8'h00;
            16'd28270: data <= 8'h1F;
            16'd28271: data <= 8'h00;
            16'd28272: data <= 8'h1F;
            16'd28273: data <= 8'h00;
            16'd28274: data <= 8'h1F;
            16'd28275: data <= 8'h00;
            16'd28276: data <= 8'h1F;
            16'd28277: data <= 8'h00;
            16'd28278: data <= 8'h1F;
            16'd28279: data <= 8'h00;
            16'd28280: data <= 8'hFF;
            16'd28281: data <= 8'hFF;
            16'd28282: data <= 8'h1F;
            16'd28283: data <= 8'h00;
            16'd28284: data <= 8'h1F;
            16'd28285: data <= 8'h00;
            16'd28286: data <= 8'h1F;
            16'd28287: data <= 8'h00;
            16'd28288: data <= 8'h1F;
            16'd28289: data <= 8'h00;
            16'd28290: data <= 8'h1F;
            16'd28291: data <= 8'h00;
            16'd28292: data <= 8'h1F;
            16'd28293: data <= 8'h00;
            16'd28294: data <= 8'h1F;
            16'd28295: data <= 8'h00;
            16'd28296: data <= 8'h1F;
            16'd28297: data <= 8'h00;
            16'd28298: data <= 8'h1F;
            16'd28299: data <= 8'h00;
            16'd28300: data <= 8'h1F;
            16'd28301: data <= 8'h00;
            16'd28302: data <= 8'h1F;
            16'd28303: data <= 8'h00;
            16'd28304: data <= 8'h1F;
            16'd28305: data <= 8'h00;
            16'd28306: data <= 8'h1F;
            16'd28307: data <= 8'h00;
            16'd28308: data <= 8'h1F;
            16'd28309: data <= 8'h00;
            16'd28310: data <= 8'h1F;
            16'd28311: data <= 8'h00;
            16'd28312: data <= 8'h1F;
            16'd28313: data <= 8'h00;
            16'd28314: data <= 8'h1F;
            16'd28315: data <= 8'h00;
            16'd28316: data <= 8'h1F;
            16'd28317: data <= 8'h00;
            16'd28318: data <= 8'h1F;
            16'd28319: data <= 8'h00;
            16'd28320: data <= 8'hFF;
            16'd28321: data <= 8'hFF;
            16'd28322: data <= 8'h1F;
            16'd28323: data <= 8'h00;
            16'd28324: data <= 8'h1F;
            16'd28325: data <= 8'h00;
            16'd28326: data <= 8'h1F;
            16'd28327: data <= 8'h00;
            16'd28328: data <= 8'h1F;
            16'd28329: data <= 8'h00;
            16'd28330: data <= 8'h1F;
            16'd28331: data <= 8'h00;
            16'd28332: data <= 8'h1F;
            16'd28333: data <= 8'h00;
            16'd28334: data <= 8'h1F;
            16'd28335: data <= 8'h00;
            16'd28336: data <= 8'h1F;
            16'd28337: data <= 8'h00;
            16'd28338: data <= 8'h1F;
            16'd28339: data <= 8'h00;
            16'd28340: data <= 8'h1F;
            16'd28341: data <= 8'h00;
            16'd28342: data <= 8'h1F;
            16'd28343: data <= 8'h00;
            16'd28344: data <= 8'h1F;
            16'd28345: data <= 8'h00;
            16'd28346: data <= 8'h1F;
            16'd28347: data <= 8'h00;
            16'd28348: data <= 8'h1F;
            16'd28349: data <= 8'h00;
            16'd28350: data <= 8'h1F;
            16'd28351: data <= 8'h00;
            16'd28352: data <= 8'h1F;
            16'd28353: data <= 8'h00;
            16'd28354: data <= 8'h1F;
            16'd28355: data <= 8'h00;
            16'd28356: data <= 8'h1F;
            16'd28357: data <= 8'h00;
            16'd28358: data <= 8'h1F;
            16'd28359: data <= 8'h00;
            16'd28360: data <= 8'hFF;
            16'd28361: data <= 8'hFF;
            16'd28362: data <= 8'h1F;
            16'd28363: data <= 8'h00;
            16'd28364: data <= 8'h1F;
            16'd28365: data <= 8'h00;
            16'd28366: data <= 8'h1F;
            16'd28367: data <= 8'h00;
            16'd28368: data <= 8'h1F;
            16'd28369: data <= 8'h00;
            16'd28370: data <= 8'h1F;
            16'd28371: data <= 8'h00;
            16'd28372: data <= 8'h1F;
            16'd28373: data <= 8'h00;
            16'd28374: data <= 8'h1F;
            16'd28375: data <= 8'h00;
            16'd28376: data <= 8'h1F;
            16'd28377: data <= 8'h00;
            16'd28378: data <= 8'h1F;
            16'd28379: data <= 8'h00;
            16'd28380: data <= 8'h1F;
            16'd28381: data <= 8'h00;
            16'd28382: data <= 8'h1F;
            16'd28383: data <= 8'h00;
            16'd28384: data <= 8'h1F;
            16'd28385: data <= 8'h00;
            16'd28386: data <= 8'h1F;
            16'd28387: data <= 8'h00;
            16'd28388: data <= 8'h1F;
            16'd28389: data <= 8'h00;
            16'd28390: data <= 8'h1F;
            16'd28391: data <= 8'h00;
            16'd28392: data <= 8'h1F;
            16'd28393: data <= 8'h00;
            16'd28394: data <= 8'h1F;
            16'd28395: data <= 8'h00;
            16'd28396: data <= 8'h1F;
            16'd28397: data <= 8'h00;
            16'd28398: data <= 8'h1F;
            16'd28399: data <= 8'h00;
            16'd28400: data <= 8'hFF;
            16'd28401: data <= 8'hFF;
            16'd28402: data <= 8'h1F;
            16'd28403: data <= 8'h00;
            16'd28404: data <= 8'h1F;
            16'd28405: data <= 8'h00;
            16'd28406: data <= 8'h1F;
            16'd28407: data <= 8'h00;
            16'd28408: data <= 8'h1F;
            16'd28409: data <= 8'h00;
            16'd28410: data <= 8'h1F;
            16'd28411: data <= 8'h00;
            16'd28412: data <= 8'h1F;
            16'd28413: data <= 8'h00;
            16'd28414: data <= 8'h1F;
            16'd28415: data <= 8'h00;
            16'd28416: data <= 8'h1F;
            16'd28417: data <= 8'h00;
            16'd28418: data <= 8'h1F;
            16'd28419: data <= 8'h00;
            16'd28420: data <= 8'h1F;
            16'd28421: data <= 8'h00;
            16'd28422: data <= 8'h1F;
            16'd28423: data <= 8'h00;
            16'd28424: data <= 8'h1F;
            16'd28425: data <= 8'h00;
            16'd28426: data <= 8'h1F;
            16'd28427: data <= 8'h00;
            16'd28428: data <= 8'h1F;
            16'd28429: data <= 8'h00;
            16'd28430: data <= 8'h1F;
            16'd28431: data <= 8'h00;
            16'd28432: data <= 8'h1F;
            16'd28433: data <= 8'h00;
            16'd28434: data <= 8'h1F;
            16'd28435: data <= 8'h00;
            16'd28436: data <= 8'h1F;
            16'd28437: data <= 8'h00;
            16'd28438: data <= 8'h1F;
            16'd28439: data <= 8'h00;
            16'd28440: data <= 8'hFF;
            16'd28441: data <= 8'hFF;
            16'd28442: data <= 8'h1F;
            16'd28443: data <= 8'h00;
            16'd28444: data <= 8'h1F;
            16'd28445: data <= 8'h00;
            16'd28446: data <= 8'h1F;
            16'd28447: data <= 8'h00;
            16'd28448: data <= 8'h1F;
            16'd28449: data <= 8'h00;
            16'd28450: data <= 8'h1F;
            16'd28451: data <= 8'h00;
            16'd28452: data <= 8'h1F;
            16'd28453: data <= 8'h00;
            16'd28454: data <= 8'h1F;
            16'd28455: data <= 8'h00;
            16'd28456: data <= 8'h1F;
            16'd28457: data <= 8'h00;
            16'd28458: data <= 8'h1F;
            16'd28459: data <= 8'h00;
            16'd28460: data <= 8'h1F;
            16'd28461: data <= 8'h00;
            16'd28462: data <= 8'h1F;
            16'd28463: data <= 8'h00;
            16'd28464: data <= 8'h1F;
            16'd28465: data <= 8'h00;
            16'd28466: data <= 8'h1F;
            16'd28467: data <= 8'h00;
            16'd28468: data <= 8'h1F;
            16'd28469: data <= 8'h00;
            16'd28470: data <= 8'h1F;
            16'd28471: data <= 8'h00;
            16'd28472: data <= 8'h1F;
            16'd28473: data <= 8'h00;
            16'd28474: data <= 8'h1F;
            16'd28475: data <= 8'h00;
            16'd28476: data <= 8'h1F;
            16'd28477: data <= 8'h00;
            16'd28478: data <= 8'h1F;
            16'd28479: data <= 8'h00;
            16'd28480: data <= 8'hFF;
            16'd28481: data <= 8'hFF;
            16'd28482: data <= 8'h1F;
            16'd28483: data <= 8'h00;
            16'd28484: data <= 8'h1F;
            16'd28485: data <= 8'h00;
            16'd28486: data <= 8'h1F;
            16'd28487: data <= 8'h00;
            16'd28488: data <= 8'h1F;
            16'd28489: data <= 8'h00;
            16'd28490: data <= 8'h1F;
            16'd28491: data <= 8'h00;
            16'd28492: data <= 8'h1F;
            16'd28493: data <= 8'h00;
            16'd28494: data <= 8'h1F;
            16'd28495: data <= 8'h00;
            16'd28496: data <= 8'h1F;
            16'd28497: data <= 8'h00;
            16'd28498: data <= 8'h1F;
            16'd28499: data <= 8'h00;
            16'd28500: data <= 8'h1F;
            16'd28501: data <= 8'h00;
            16'd28502: data <= 8'h1F;
            16'd28503: data <= 8'h00;
            16'd28504: data <= 8'h1F;
            16'd28505: data <= 8'h00;
            16'd28506: data <= 8'h1F;
            16'd28507: data <= 8'h00;
            16'd28508: data <= 8'h1F;
            16'd28509: data <= 8'h00;
            16'd28510: data <= 8'h1F;
            16'd28511: data <= 8'h00;
            16'd28512: data <= 8'h1F;
            16'd28513: data <= 8'h00;
            16'd28514: data <= 8'h1F;
            16'd28515: data <= 8'h00;
            16'd28516: data <= 8'h1F;
            16'd28517: data <= 8'h00;
            16'd28518: data <= 8'h1F;
            16'd28519: data <= 8'h00;
            16'd28520: data <= 8'hFF;
            16'd28521: data <= 8'hFF;
            16'd28522: data <= 8'h1F;
            16'd28523: data <= 8'h00;
            16'd28524: data <= 8'h1F;
            16'd28525: data <= 8'h00;
            16'd28526: data <= 8'h1F;
            16'd28527: data <= 8'h00;
            16'd28528: data <= 8'h1F;
            16'd28529: data <= 8'h00;
            16'd28530: data <= 8'h1F;
            16'd28531: data <= 8'h00;
            16'd28532: data <= 8'h1F;
            16'd28533: data <= 8'h00;
            16'd28534: data <= 8'h1F;
            16'd28535: data <= 8'h00;
            16'd28536: data <= 8'h1F;
            16'd28537: data <= 8'h00;
            16'd28538: data <= 8'h1F;
            16'd28539: data <= 8'h00;
            16'd28540: data <= 8'h1F;
            16'd28541: data <= 8'h00;
            16'd28542: data <= 8'h1F;
            16'd28543: data <= 8'h00;
            16'd28544: data <= 8'h1F;
            16'd28545: data <= 8'h00;
            16'd28546: data <= 8'h1F;
            16'd28547: data <= 8'h00;
            16'd28548: data <= 8'h1F;
            16'd28549: data <= 8'h00;
            16'd28550: data <= 8'h1F;
            16'd28551: data <= 8'h00;
            16'd28552: data <= 8'h1F;
            16'd28553: data <= 8'h00;
            16'd28554: data <= 8'h1F;
            16'd28555: data <= 8'h00;
            16'd28556: data <= 8'h1F;
            16'd28557: data <= 8'h00;
            16'd28558: data <= 8'h1F;
            16'd28559: data <= 8'h00;
            16'd28560: data <= 8'hFF;
            16'd28561: data <= 8'hFF;
            16'd28562: data <= 8'h1F;
            16'd28563: data <= 8'h00;
            16'd28564: data <= 8'h1F;
            16'd28565: data <= 8'h00;
            16'd28566: data <= 8'h1F;
            16'd28567: data <= 8'h00;
            16'd28568: data <= 8'h1F;
            16'd28569: data <= 8'h00;
            16'd28570: data <= 8'h1F;
            16'd28571: data <= 8'h00;
            16'd28572: data <= 8'h1F;
            16'd28573: data <= 8'h00;
            16'd28574: data <= 8'h1F;
            16'd28575: data <= 8'h00;
            16'd28576: data <= 8'h1F;
            16'd28577: data <= 8'h00;
            16'd28578: data <= 8'h1F;
            16'd28579: data <= 8'h00;
            16'd28580: data <= 8'h1F;
            16'd28581: data <= 8'h00;
            16'd28582: data <= 8'h1F;
            16'd28583: data <= 8'h00;
            16'd28584: data <= 8'h1F;
            16'd28585: data <= 8'h00;
            16'd28586: data <= 8'h1F;
            16'd28587: data <= 8'h00;
            16'd28588: data <= 8'h1F;
            16'd28589: data <= 8'h00;
            16'd28590: data <= 8'h1F;
            16'd28591: data <= 8'h00;
            16'd28592: data <= 8'h1F;
            16'd28593: data <= 8'h00;
            16'd28594: data <= 8'h1F;
            16'd28595: data <= 8'h00;
            16'd28596: data <= 8'h1F;
            16'd28597: data <= 8'h00;
            16'd28598: data <= 8'h1F;
            16'd28599: data <= 8'h00;
            16'd28600: data <= 8'hFF;
            16'd28601: data <= 8'hFF;
            16'd28602: data <= 8'h1F;
            16'd28603: data <= 8'h00;
            16'd28604: data <= 8'h1F;
            16'd28605: data <= 8'h00;
            16'd28606: data <= 8'h1F;
            16'd28607: data <= 8'h00;
            16'd28608: data <= 8'h1F;
            16'd28609: data <= 8'h00;
            16'd28610: data <= 8'h1F;
            16'd28611: data <= 8'h00;
            16'd28612: data <= 8'h1F;
            16'd28613: data <= 8'h00;
            16'd28614: data <= 8'h1F;
            16'd28615: data <= 8'h00;
            16'd28616: data <= 8'h1F;
            16'd28617: data <= 8'h00;
            16'd28618: data <= 8'h1F;
            16'd28619: data <= 8'h00;
            16'd28620: data <= 8'h1F;
            16'd28621: data <= 8'h00;
            16'd28622: data <= 8'h1F;
            16'd28623: data <= 8'h00;
            16'd28624: data <= 8'h1F;
            16'd28625: data <= 8'h00;
            16'd28626: data <= 8'h1F;
            16'd28627: data <= 8'h00;
            16'd28628: data <= 8'h1F;
            16'd28629: data <= 8'h00;
            16'd28630: data <= 8'h1F;
            16'd28631: data <= 8'h00;
            16'd28632: data <= 8'h1F;
            16'd28633: data <= 8'h00;
            16'd28634: data <= 8'h1F;
            16'd28635: data <= 8'h00;
            16'd28636: data <= 8'h1F;
            16'd28637: data <= 8'h00;
            16'd28638: data <= 8'h1F;
            16'd28639: data <= 8'h00;
            16'd28640: data <= 8'hFF;
            16'd28641: data <= 8'hFF;
            16'd28642: data <= 8'h1F;
            16'd28643: data <= 8'h00;
            16'd28644: data <= 8'h1F;
            16'd28645: data <= 8'h00;
            16'd28646: data <= 8'h1F;
            16'd28647: data <= 8'h00;
            16'd28648: data <= 8'h1F;
            16'd28649: data <= 8'h00;
            16'd28650: data <= 8'h1F;
            16'd28651: data <= 8'h00;
            16'd28652: data <= 8'h1F;
            16'd28653: data <= 8'h00;
            16'd28654: data <= 8'h1F;
            16'd28655: data <= 8'h00;
            16'd28656: data <= 8'h1F;
            16'd28657: data <= 8'h00;
            16'd28658: data <= 8'h1F;
            16'd28659: data <= 8'h00;
            16'd28660: data <= 8'h1F;
            16'd28661: data <= 8'h00;
            16'd28662: data <= 8'h1F;
            16'd28663: data <= 8'h00;
            16'd28664: data <= 8'h1F;
            16'd28665: data <= 8'h00;
            16'd28666: data <= 8'h1F;
            16'd28667: data <= 8'h00;
            16'd28668: data <= 8'h1F;
            16'd28669: data <= 8'h00;
            16'd28670: data <= 8'h1F;
            16'd28671: data <= 8'h00;
            16'd28672: data <= 8'h1F;
            16'd28673: data <= 8'h00;
            16'd28674: data <= 8'h1F;
            16'd28675: data <= 8'h00;
            16'd28676: data <= 8'h1F;
            16'd28677: data <= 8'h00;
            16'd28678: data <= 8'h1F;
            16'd28679: data <= 8'h00;
            16'd28680: data <= 8'hFF;
            16'd28681: data <= 8'hFF;
            16'd28682: data <= 8'h1F;
            16'd28683: data <= 8'h00;
            16'd28684: data <= 8'h1F;
            16'd28685: data <= 8'h00;
            16'd28686: data <= 8'h1F;
            16'd28687: data <= 8'h00;
            16'd28688: data <= 8'h1F;
            16'd28689: data <= 8'h00;
            16'd28690: data <= 8'h1F;
            16'd28691: data <= 8'h00;
            16'd28692: data <= 8'h1F;
            16'd28693: data <= 8'h00;
            16'd28694: data <= 8'h1F;
            16'd28695: data <= 8'h00;
            16'd28696: data <= 8'h1F;
            16'd28697: data <= 8'h00;
            16'd28698: data <= 8'h1F;
            16'd28699: data <= 8'h00;
            16'd28700: data <= 8'h1F;
            16'd28701: data <= 8'h00;
            16'd28702: data <= 8'h1F;
            16'd28703: data <= 8'h00;
            16'd28704: data <= 8'h1F;
            16'd28705: data <= 8'h00;
            16'd28706: data <= 8'h1F;
            16'd28707: data <= 8'h00;
            16'd28708: data <= 8'h1F;
            16'd28709: data <= 8'h00;
            16'd28710: data <= 8'h1F;
            16'd28711: data <= 8'h00;
            16'd28712: data <= 8'h1F;
            16'd28713: data <= 8'h00;
            16'd28714: data <= 8'h1F;
            16'd28715: data <= 8'h00;
            16'd28716: data <= 8'h1F;
            16'd28717: data <= 8'h00;
            16'd28718: data <= 8'h1F;
            16'd28719: data <= 8'h00;
            16'd28720: data <= 8'hFF;
            16'd28721: data <= 8'hFF;
            16'd28722: data <= 8'h1F;
            16'd28723: data <= 8'h00;
            16'd28724: data <= 8'h1F;
            16'd28725: data <= 8'h00;
            16'd28726: data <= 8'h1F;
            16'd28727: data <= 8'h00;
            16'd28728: data <= 8'h1F;
            16'd28729: data <= 8'h00;
            16'd28730: data <= 8'h1F;
            16'd28731: data <= 8'h00;
            16'd28732: data <= 8'h1F;
            16'd28733: data <= 8'h00;
            16'd28734: data <= 8'h1F;
            16'd28735: data <= 8'h00;
            16'd28736: data <= 8'h1F;
            16'd28737: data <= 8'h00;
            16'd28738: data <= 8'h1F;
            16'd28739: data <= 8'h00;
            16'd28740: data <= 8'h1F;
            16'd28741: data <= 8'h00;
            16'd28742: data <= 8'h1F;
            16'd28743: data <= 8'h00;
            16'd28744: data <= 8'h1F;
            16'd28745: data <= 8'h00;
            16'd28746: data <= 8'h1F;
            16'd28747: data <= 8'h00;
            16'd28748: data <= 8'h1F;
            16'd28749: data <= 8'h00;
            16'd28750: data <= 8'h1F;
            16'd28751: data <= 8'h00;
            16'd28752: data <= 8'h1F;
            16'd28753: data <= 8'h00;
            16'd28754: data <= 8'h1F;
            16'd28755: data <= 8'h00;
            16'd28756: data <= 8'h1F;
            16'd28757: data <= 8'h00;
            16'd28758: data <= 8'h1F;
            16'd28759: data <= 8'h00;
            16'd28760: data <= 8'hFF;
            16'd28761: data <= 8'hFF;
            16'd28762: data <= 8'h1F;
            16'd28763: data <= 8'h00;
            16'd28764: data <= 8'h1F;
            16'd28765: data <= 8'h00;
            16'd28766: data <= 8'h1F;
            16'd28767: data <= 8'h00;
            16'd28768: data <= 8'h1F;
            16'd28769: data <= 8'h00;
            16'd28770: data <= 8'h1F;
            16'd28771: data <= 8'h00;
            16'd28772: data <= 8'h1F;
            16'd28773: data <= 8'h00;
            16'd28774: data <= 8'h1F;
            16'd28775: data <= 8'h00;
            16'd28776: data <= 8'h1F;
            16'd28777: data <= 8'h00;
            16'd28778: data <= 8'h1F;
            16'd28779: data <= 8'h00;
            16'd28780: data <= 8'h1F;
            16'd28781: data <= 8'h00;
            16'd28782: data <= 8'h1F;
            16'd28783: data <= 8'h00;
            16'd28784: data <= 8'h1F;
            16'd28785: data <= 8'h00;
            16'd28786: data <= 8'h1F;
            16'd28787: data <= 8'h00;
            16'd28788: data <= 8'h1F;
            16'd28789: data <= 8'h00;
            16'd28790: data <= 8'h1F;
            16'd28791: data <= 8'h00;
            16'd28792: data <= 8'h1F;
            16'd28793: data <= 8'h00;
            16'd28794: data <= 8'h1F;
            16'd28795: data <= 8'h00;
            16'd28796: data <= 8'h1F;
            16'd28797: data <= 8'h00;
            16'd28798: data <= 8'h1F;
            16'd28799: data <= 8'h00;
            16'd28800: data <= 8'hFF;
            16'd28801: data <= 8'hFF;
            16'd28802: data <= 8'hFF;
            16'd28803: data <= 8'hFF;
            16'd28804: data <= 8'hFF;
            16'd28805: data <= 8'hFF;
            16'd28806: data <= 8'hFF;
            16'd28807: data <= 8'hFF;
            16'd28808: data <= 8'hFF;
            16'd28809: data <= 8'hFF;
            16'd28810: data <= 8'hFF;
            16'd28811: data <= 8'hFF;
            16'd28812: data <= 8'hFF;
            16'd28813: data <= 8'hFF;
            16'd28814: data <= 8'hFF;
            16'd28815: data <= 8'hFF;
            16'd28816: data <= 8'hFF;
            16'd28817: data <= 8'hFF;
            16'd28818: data <= 8'hFF;
            16'd28819: data <= 8'hFF;
            16'd28820: data <= 8'hFF;
            16'd28821: data <= 8'hFF;
            16'd28822: data <= 8'hFF;
            16'd28823: data <= 8'hFF;
            16'd28824: data <= 8'hFF;
            16'd28825: data <= 8'hFF;
            16'd28826: data <= 8'hFF;
            16'd28827: data <= 8'hFF;
            16'd28828: data <= 8'hFF;
            16'd28829: data <= 8'hFF;
            16'd28830: data <= 8'hFF;
            16'd28831: data <= 8'hFF;
            16'd28832: data <= 8'hFF;
            16'd28833: data <= 8'hFF;
            16'd28834: data <= 8'hFF;
            16'd28835: data <= 8'hFF;
            16'd28836: data <= 8'hFF;
            16'd28837: data <= 8'hFF;
            16'd28838: data <= 8'hFF;
            16'd28839: data <= 8'hFF;
            16'd28840: data <= 8'hFF;
            16'd28841: data <= 8'hFF;
            16'd28842: data <= 8'hFF;
            16'd28843: data <= 8'hFF;
            16'd28844: data <= 8'hFF;
            16'd28845: data <= 8'hFF;
            16'd28846: data <= 8'hFF;
            16'd28847: data <= 8'hFF;
            16'd28848: data <= 8'hFF;
            16'd28849: data <= 8'hFF;
            16'd28850: data <= 8'hFF;
            16'd28851: data <= 8'hFF;
            16'd28852: data <= 8'hFF;
            16'd28853: data <= 8'hFF;
            16'd28854: data <= 8'hFF;
            16'd28855: data <= 8'hFF;
            16'd28856: data <= 8'hFF;
            16'd28857: data <= 8'hFF;
            16'd28858: data <= 8'hFF;
            16'd28859: data <= 8'hFF;
            16'd28860: data <= 8'hFF;
            16'd28861: data <= 8'hFF;
            16'd28862: data <= 8'hFF;
            16'd28863: data <= 8'hFF;
            16'd28864: data <= 8'hFF;
            16'd28865: data <= 8'hFF;
            16'd28866: data <= 8'hFF;
            16'd28867: data <= 8'hFF;
            16'd28868: data <= 8'hFF;
            16'd28869: data <= 8'hFF;
            16'd28870: data <= 8'hFF;
            16'd28871: data <= 8'hFF;
            16'd28872: data <= 8'hFF;
            16'd28873: data <= 8'hFF;
            16'd28874: data <= 8'hFF;
            16'd28875: data <= 8'hFF;
            16'd28876: data <= 8'hFF;
            16'd28877: data <= 8'hFF;
            16'd28878: data <= 8'hFF;
            16'd28879: data <= 8'hFF;
            16'd28880: data <= 8'hFF;
            16'd28881: data <= 8'hFF;
            16'd28882: data <= 8'hFF;
            16'd28883: data <= 8'hFF;
            16'd28884: data <= 8'hFF;
            16'd28885: data <= 8'hFF;
            16'd28886: data <= 8'hFF;
            16'd28887: data <= 8'hFF;
            16'd28888: data <= 8'hFF;
            16'd28889: data <= 8'hFF;
            16'd28890: data <= 8'hFF;
            16'd28891: data <= 8'hFF;
            16'd28892: data <= 8'hFF;
            16'd28893: data <= 8'hFF;
            16'd28894: data <= 8'hFF;
            16'd28895: data <= 8'hFF;
            16'd28896: data <= 8'hFF;
            16'd28897: data <= 8'hFF;
            16'd28898: data <= 8'hFF;
            16'd28899: data <= 8'hFF;
            16'd28900: data <= 8'hFF;
            16'd28901: data <= 8'hFF;
            16'd28902: data <= 8'hFF;
            16'd28903: data <= 8'hFF;
            16'd28904: data <= 8'hFF;
            16'd28905: data <= 8'hFF;
            16'd28906: data <= 8'hFF;
            16'd28907: data <= 8'hFF;
            16'd28908: data <= 8'hFF;
            16'd28909: data <= 8'hFF;
            16'd28910: data <= 8'hFF;
            16'd28911: data <= 8'hFF;
            16'd28912: data <= 8'hFF;
            16'd28913: data <= 8'hFF;
            16'd28914: data <= 8'hFF;
            16'd28915: data <= 8'hFF;
            16'd28916: data <= 8'hFF;
            16'd28917: data <= 8'hFF;
            16'd28918: data <= 8'hFF;
            16'd28919: data <= 8'hFF;
            16'd28920: data <= 8'hFF;
            16'd28921: data <= 8'hFF;
            16'd28922: data <= 8'hFF;
            16'd28923: data <= 8'hFF;
            16'd28924: data <= 8'hFF;
            16'd28925: data <= 8'hFF;
            16'd28926: data <= 8'hFF;
            16'd28927: data <= 8'hFF;
            16'd28928: data <= 8'hFF;
            16'd28929: data <= 8'hFF;
            16'd28930: data <= 8'hFF;
            16'd28931: data <= 8'hFF;
            16'd28932: data <= 8'hFF;
            16'd28933: data <= 8'hFF;
            16'd28934: data <= 8'hFF;
            16'd28935: data <= 8'hFF;
            16'd28936: data <= 8'hFF;
            16'd28937: data <= 8'hFF;
            16'd28938: data <= 8'hFF;
            16'd28939: data <= 8'hFF;
            16'd28940: data <= 8'hFF;
            16'd28941: data <= 8'hFF;
            16'd28942: data <= 8'hFF;
            16'd28943: data <= 8'hFF;
            16'd28944: data <= 8'hFF;
            16'd28945: data <= 8'hFF;
            16'd28946: data <= 8'hFF;
            16'd28947: data <= 8'hFF;
            16'd28948: data <= 8'hFF;
            16'd28949: data <= 8'hFF;
            16'd28950: data <= 8'hFF;
            16'd28951: data <= 8'hFF;
            16'd28952: data <= 8'hFF;
            16'd28953: data <= 8'hFF;
            16'd28954: data <= 8'hFF;
            16'd28955: data <= 8'hFF;
            16'd28956: data <= 8'hFF;
            16'd28957: data <= 8'hFF;
            16'd28958: data <= 8'hFF;
            16'd28959: data <= 8'hFF;
            16'd28960: data <= 8'hFF;
            16'd28961: data <= 8'hFF;
            16'd28962: data <= 8'hFF;
            16'd28963: data <= 8'hFF;
            16'd28964: data <= 8'hFF;
            16'd28965: data <= 8'hFF;
            16'd28966: data <= 8'hFF;
            16'd28967: data <= 8'hFF;
            16'd28968: data <= 8'hFF;
            16'd28969: data <= 8'hFF;
            16'd28970: data <= 8'hFF;
            16'd28971: data <= 8'hFF;
            16'd28972: data <= 8'hFF;
            16'd28973: data <= 8'hFF;
            16'd28974: data <= 8'hFF;
            16'd28975: data <= 8'hFF;
            16'd28976: data <= 8'hFF;
            16'd28977: data <= 8'hFF;
            16'd28978: data <= 8'hFF;
            16'd28979: data <= 8'hFF;
            16'd28980: data <= 8'hFF;
            16'd28981: data <= 8'hFF;
            16'd28982: data <= 8'hFF;
            16'd28983: data <= 8'hFF;
            16'd28984: data <= 8'hFF;
            16'd28985: data <= 8'hFF;
            16'd28986: data <= 8'hFF;
            16'd28987: data <= 8'hFF;
            16'd28988: data <= 8'hFF;
            16'd28989: data <= 8'hFF;
            16'd28990: data <= 8'hFF;
            16'd28991: data <= 8'hFF;
            16'd28992: data <= 8'hFF;
            16'd28993: data <= 8'hFF;
            16'd28994: data <= 8'hFF;
            16'd28995: data <= 8'hFF;
            16'd28996: data <= 8'hFF;
            16'd28997: data <= 8'hFF;
            16'd28998: data <= 8'hFF;
            16'd28999: data <= 8'hFF;
            16'd29000: data <= 8'hFF;
            16'd29001: data <= 8'hFF;
            16'd29002: data <= 8'hFF;
            16'd29003: data <= 8'hFF;
            16'd29004: data <= 8'hFF;
            16'd29005: data <= 8'hFF;
            16'd29006: data <= 8'hFF;
            16'd29007: data <= 8'hFF;
            16'd29008: data <= 8'hFF;
            16'd29009: data <= 8'hFF;
            16'd29010: data <= 8'hFF;
            16'd29011: data <= 8'hFF;
            16'd29012: data <= 8'hFF;
            16'd29013: data <= 8'hFF;
            16'd29014: data <= 8'hFF;
            16'd29015: data <= 8'hFF;
            16'd29016: data <= 8'hFF;
            16'd29017: data <= 8'hFF;
            16'd29018: data <= 8'hFF;
            16'd29019: data <= 8'hFF;
            16'd29020: data <= 8'hFF;
            16'd29021: data <= 8'hFF;
            16'd29022: data <= 8'hFF;
            16'd29023: data <= 8'hFF;
            16'd29024: data <= 8'hFF;
            16'd29025: data <= 8'hFF;
            16'd29026: data <= 8'hFF;
            16'd29027: data <= 8'hFF;
            16'd29028: data <= 8'hFF;
            16'd29029: data <= 8'hFF;
            16'd29030: data <= 8'hFF;
            16'd29031: data <= 8'hFF;
            16'd29032: data <= 8'hFF;
            16'd29033: data <= 8'hFF;
            16'd29034: data <= 8'hFF;
            16'd29035: data <= 8'hFF;
            16'd29036: data <= 8'hFF;
            16'd29037: data <= 8'hFF;
            16'd29038: data <= 8'hFF;
            16'd29039: data <= 8'hFF;
            16'd29040: data <= 8'hFF;
            16'd29041: data <= 8'hFF;
            16'd29042: data <= 8'h1F;
            16'd29043: data <= 8'h00;
            16'd29044: data <= 8'h1F;
            16'd29045: data <= 8'h00;
            16'd29046: data <= 8'h1F;
            16'd29047: data <= 8'h00;
            16'd29048: data <= 8'h1F;
            16'd29049: data <= 8'h00;
            16'd29050: data <= 8'h1F;
            16'd29051: data <= 8'h00;
            16'd29052: data <= 8'h1F;
            16'd29053: data <= 8'h00;
            16'd29054: data <= 8'h1F;
            16'd29055: data <= 8'h00;
            16'd29056: data <= 8'h1F;
            16'd29057: data <= 8'h00;
            16'd29058: data <= 8'h1F;
            16'd29059: data <= 8'h00;
            16'd29060: data <= 8'h1F;
            16'd29061: data <= 8'h00;
            16'd29062: data <= 8'h1F;
            16'd29063: data <= 8'h00;
            16'd29064: data <= 8'h1F;
            16'd29065: data <= 8'h00;
            16'd29066: data <= 8'h1F;
            16'd29067: data <= 8'h00;
            16'd29068: data <= 8'h1F;
            16'd29069: data <= 8'h00;
            16'd29070: data <= 8'h1F;
            16'd29071: data <= 8'h00;
            16'd29072: data <= 8'h1F;
            16'd29073: data <= 8'h00;
            16'd29074: data <= 8'h1F;
            16'd29075: data <= 8'h00;
            16'd29076: data <= 8'h1F;
            16'd29077: data <= 8'h00;
            16'd29078: data <= 8'h1F;
            16'd29079: data <= 8'h00;
            16'd29080: data <= 8'hFF;
            16'd29081: data <= 8'hFF;
            16'd29082: data <= 8'h1F;
            16'd29083: data <= 8'h00;
            16'd29084: data <= 8'h1F;
            16'd29085: data <= 8'h00;
            16'd29086: data <= 8'h1F;
            16'd29087: data <= 8'h00;
            16'd29088: data <= 8'h1F;
            16'd29089: data <= 8'h00;
            16'd29090: data <= 8'h1F;
            16'd29091: data <= 8'h00;
            16'd29092: data <= 8'h1F;
            16'd29093: data <= 8'h00;
            16'd29094: data <= 8'h1F;
            16'd29095: data <= 8'h00;
            16'd29096: data <= 8'h1F;
            16'd29097: data <= 8'h00;
            16'd29098: data <= 8'h1F;
            16'd29099: data <= 8'h00;
            16'd29100: data <= 8'h1F;
            16'd29101: data <= 8'h00;
            16'd29102: data <= 8'h1F;
            16'd29103: data <= 8'h00;
            16'd29104: data <= 8'h1F;
            16'd29105: data <= 8'h00;
            16'd29106: data <= 8'h1F;
            16'd29107: data <= 8'h00;
            16'd29108: data <= 8'h1F;
            16'd29109: data <= 8'h00;
            16'd29110: data <= 8'h1F;
            16'd29111: data <= 8'h00;
            16'd29112: data <= 8'h1F;
            16'd29113: data <= 8'h00;
            16'd29114: data <= 8'h1F;
            16'd29115: data <= 8'h00;
            16'd29116: data <= 8'h1F;
            16'd29117: data <= 8'h00;
            16'd29118: data <= 8'h1F;
            16'd29119: data <= 8'h00;
            16'd29120: data <= 8'hFF;
            16'd29121: data <= 8'hFF;
            16'd29122: data <= 8'h1F;
            16'd29123: data <= 8'h00;
            16'd29124: data <= 8'h1F;
            16'd29125: data <= 8'h00;
            16'd29126: data <= 8'h1F;
            16'd29127: data <= 8'h00;
            16'd29128: data <= 8'h1F;
            16'd29129: data <= 8'h00;
            16'd29130: data <= 8'h1F;
            16'd29131: data <= 8'h00;
            16'd29132: data <= 8'h1F;
            16'd29133: data <= 8'h00;
            16'd29134: data <= 8'h1F;
            16'd29135: data <= 8'h00;
            16'd29136: data <= 8'h1F;
            16'd29137: data <= 8'h00;
            16'd29138: data <= 8'h1F;
            16'd29139: data <= 8'h00;
            16'd29140: data <= 8'h1F;
            16'd29141: data <= 8'h00;
            16'd29142: data <= 8'h1F;
            16'd29143: data <= 8'h00;
            16'd29144: data <= 8'h1F;
            16'd29145: data <= 8'h00;
            16'd29146: data <= 8'h1F;
            16'd29147: data <= 8'h00;
            16'd29148: data <= 8'h1F;
            16'd29149: data <= 8'h00;
            16'd29150: data <= 8'h1F;
            16'd29151: data <= 8'h00;
            16'd29152: data <= 8'h1F;
            16'd29153: data <= 8'h00;
            16'd29154: data <= 8'h1F;
            16'd29155: data <= 8'h00;
            16'd29156: data <= 8'h1F;
            16'd29157: data <= 8'h00;
            16'd29158: data <= 8'h1F;
            16'd29159: data <= 8'h00;
            16'd29160: data <= 8'hFF;
            16'd29161: data <= 8'hFF;
            16'd29162: data <= 8'h1F;
            16'd29163: data <= 8'h00;
            16'd29164: data <= 8'h1F;
            16'd29165: data <= 8'h00;
            16'd29166: data <= 8'h1F;
            16'd29167: data <= 8'h00;
            16'd29168: data <= 8'h1F;
            16'd29169: data <= 8'h00;
            16'd29170: data <= 8'h1F;
            16'd29171: data <= 8'h00;
            16'd29172: data <= 8'h1F;
            16'd29173: data <= 8'h00;
            16'd29174: data <= 8'h1F;
            16'd29175: data <= 8'h00;
            16'd29176: data <= 8'h1F;
            16'd29177: data <= 8'h00;
            16'd29178: data <= 8'h1F;
            16'd29179: data <= 8'h00;
            16'd29180: data <= 8'h1F;
            16'd29181: data <= 8'h00;
            16'd29182: data <= 8'h1F;
            16'd29183: data <= 8'h00;
            16'd29184: data <= 8'h1F;
            16'd29185: data <= 8'h00;
            16'd29186: data <= 8'h1F;
            16'd29187: data <= 8'h00;
            16'd29188: data <= 8'h1F;
            16'd29189: data <= 8'h00;
            16'd29190: data <= 8'h1F;
            16'd29191: data <= 8'h00;
            16'd29192: data <= 8'h1F;
            16'd29193: data <= 8'h00;
            16'd29194: data <= 8'h1F;
            16'd29195: data <= 8'h00;
            16'd29196: data <= 8'h1F;
            16'd29197: data <= 8'h00;
            16'd29198: data <= 8'h1F;
            16'd29199: data <= 8'h00;
            16'd29200: data <= 8'hFF;
            16'd29201: data <= 8'hFF;
            16'd29202: data <= 8'h1F;
            16'd29203: data <= 8'h00;
            16'd29204: data <= 8'h1F;
            16'd29205: data <= 8'h00;
            16'd29206: data <= 8'h1F;
            16'd29207: data <= 8'h00;
            16'd29208: data <= 8'h1F;
            16'd29209: data <= 8'h00;
            16'd29210: data <= 8'h1F;
            16'd29211: data <= 8'h00;
            16'd29212: data <= 8'h1F;
            16'd29213: data <= 8'h00;
            16'd29214: data <= 8'h1F;
            16'd29215: data <= 8'h00;
            16'd29216: data <= 8'h1F;
            16'd29217: data <= 8'h00;
            16'd29218: data <= 8'h1F;
            16'd29219: data <= 8'h00;
            16'd29220: data <= 8'h1F;
            16'd29221: data <= 8'h00;
            16'd29222: data <= 8'h1F;
            16'd29223: data <= 8'h00;
            16'd29224: data <= 8'h1F;
            16'd29225: data <= 8'h00;
            16'd29226: data <= 8'h1F;
            16'd29227: data <= 8'h00;
            16'd29228: data <= 8'h1F;
            16'd29229: data <= 8'h00;
            16'd29230: data <= 8'h1F;
            16'd29231: data <= 8'h00;
            16'd29232: data <= 8'h1F;
            16'd29233: data <= 8'h00;
            16'd29234: data <= 8'h1F;
            16'd29235: data <= 8'h00;
            16'd29236: data <= 8'h1F;
            16'd29237: data <= 8'h00;
            16'd29238: data <= 8'h1F;
            16'd29239: data <= 8'h00;
            16'd29240: data <= 8'hFF;
            16'd29241: data <= 8'hFF;
            16'd29242: data <= 8'h1F;
            16'd29243: data <= 8'h00;
            16'd29244: data <= 8'h1F;
            16'd29245: data <= 8'h00;
            16'd29246: data <= 8'h1F;
            16'd29247: data <= 8'h00;
            16'd29248: data <= 8'h1F;
            16'd29249: data <= 8'h00;
            16'd29250: data <= 8'h1F;
            16'd29251: data <= 8'h00;
            16'd29252: data <= 8'h1F;
            16'd29253: data <= 8'h00;
            16'd29254: data <= 8'h1F;
            16'd29255: data <= 8'h00;
            16'd29256: data <= 8'h1F;
            16'd29257: data <= 8'h00;
            16'd29258: data <= 8'h1F;
            16'd29259: data <= 8'h00;
            16'd29260: data <= 8'h1F;
            16'd29261: data <= 8'h00;
            16'd29262: data <= 8'h1F;
            16'd29263: data <= 8'h00;
            16'd29264: data <= 8'h1F;
            16'd29265: data <= 8'h00;
            16'd29266: data <= 8'h1F;
            16'd29267: data <= 8'h00;
            16'd29268: data <= 8'h1F;
            16'd29269: data <= 8'h00;
            16'd29270: data <= 8'h1F;
            16'd29271: data <= 8'h00;
            16'd29272: data <= 8'h1F;
            16'd29273: data <= 8'h00;
            16'd29274: data <= 8'h1F;
            16'd29275: data <= 8'h00;
            16'd29276: data <= 8'h1F;
            16'd29277: data <= 8'h00;
            16'd29278: data <= 8'h1F;
            16'd29279: data <= 8'h00;
            16'd29280: data <= 8'hFF;
            16'd29281: data <= 8'hFF;
            16'd29282: data <= 8'h1F;
            16'd29283: data <= 8'h00;
            16'd29284: data <= 8'h1F;
            16'd29285: data <= 8'h00;
            16'd29286: data <= 8'h1F;
            16'd29287: data <= 8'h00;
            16'd29288: data <= 8'h1F;
            16'd29289: data <= 8'h00;
            16'd29290: data <= 8'h1F;
            16'd29291: data <= 8'h00;
            16'd29292: data <= 8'h1F;
            16'd29293: data <= 8'h00;
            16'd29294: data <= 8'h1F;
            16'd29295: data <= 8'h00;
            16'd29296: data <= 8'h1F;
            16'd29297: data <= 8'h00;
            16'd29298: data <= 8'h1F;
            16'd29299: data <= 8'h00;
            16'd29300: data <= 8'h1F;
            16'd29301: data <= 8'h00;
            16'd29302: data <= 8'h1F;
            16'd29303: data <= 8'h00;
            16'd29304: data <= 8'h1F;
            16'd29305: data <= 8'h00;
            16'd29306: data <= 8'h1F;
            16'd29307: data <= 8'h00;
            16'd29308: data <= 8'h1F;
            16'd29309: data <= 8'h00;
            16'd29310: data <= 8'h1F;
            16'd29311: data <= 8'h00;
            16'd29312: data <= 8'h1F;
            16'd29313: data <= 8'h00;
            16'd29314: data <= 8'h1F;
            16'd29315: data <= 8'h00;
            16'd29316: data <= 8'h1F;
            16'd29317: data <= 8'h00;
            16'd29318: data <= 8'h1F;
            16'd29319: data <= 8'h00;
            16'd29320: data <= 8'hFF;
            16'd29321: data <= 8'hFF;
            16'd29322: data <= 8'h1F;
            16'd29323: data <= 8'h00;
            16'd29324: data <= 8'h1F;
            16'd29325: data <= 8'h00;
            16'd29326: data <= 8'h1F;
            16'd29327: data <= 8'h00;
            16'd29328: data <= 8'h1F;
            16'd29329: data <= 8'h00;
            16'd29330: data <= 8'h1F;
            16'd29331: data <= 8'h00;
            16'd29332: data <= 8'h1F;
            16'd29333: data <= 8'h00;
            16'd29334: data <= 8'h1F;
            16'd29335: data <= 8'h00;
            16'd29336: data <= 8'h1F;
            16'd29337: data <= 8'h00;
            16'd29338: data <= 8'h1F;
            16'd29339: data <= 8'h00;
            16'd29340: data <= 8'h1F;
            16'd29341: data <= 8'h00;
            16'd29342: data <= 8'h1F;
            16'd29343: data <= 8'h00;
            16'd29344: data <= 8'h1F;
            16'd29345: data <= 8'h00;
            16'd29346: data <= 8'h1F;
            16'd29347: data <= 8'h00;
            16'd29348: data <= 8'h1F;
            16'd29349: data <= 8'h00;
            16'd29350: data <= 8'h1F;
            16'd29351: data <= 8'h00;
            16'd29352: data <= 8'h1F;
            16'd29353: data <= 8'h00;
            16'd29354: data <= 8'h1F;
            16'd29355: data <= 8'h00;
            16'd29356: data <= 8'h1F;
            16'd29357: data <= 8'h00;
            16'd29358: data <= 8'h1F;
            16'd29359: data <= 8'h00;
            16'd29360: data <= 8'hFF;
            16'd29361: data <= 8'hFF;
            16'd29362: data <= 8'h1F;
            16'd29363: data <= 8'h00;
            16'd29364: data <= 8'h1F;
            16'd29365: data <= 8'h00;
            16'd29366: data <= 8'h1F;
            16'd29367: data <= 8'h00;
            16'd29368: data <= 8'h1F;
            16'd29369: data <= 8'h00;
            16'd29370: data <= 8'h1F;
            16'd29371: data <= 8'h00;
            16'd29372: data <= 8'h1F;
            16'd29373: data <= 8'h00;
            16'd29374: data <= 8'h1F;
            16'd29375: data <= 8'h00;
            16'd29376: data <= 8'h1F;
            16'd29377: data <= 8'h00;
            16'd29378: data <= 8'h1F;
            16'd29379: data <= 8'h00;
            16'd29380: data <= 8'h1F;
            16'd29381: data <= 8'h00;
            16'd29382: data <= 8'h1F;
            16'd29383: data <= 8'h00;
            16'd29384: data <= 8'h1F;
            16'd29385: data <= 8'h00;
            16'd29386: data <= 8'h1F;
            16'd29387: data <= 8'h00;
            16'd29388: data <= 8'h1F;
            16'd29389: data <= 8'h00;
            16'd29390: data <= 8'h1F;
            16'd29391: data <= 8'h00;
            16'd29392: data <= 8'h1F;
            16'd29393: data <= 8'h00;
            16'd29394: data <= 8'h1F;
            16'd29395: data <= 8'h00;
            16'd29396: data <= 8'h1F;
            16'd29397: data <= 8'h00;
            16'd29398: data <= 8'h1F;
            16'd29399: data <= 8'h00;
            16'd29400: data <= 8'hFF;
            16'd29401: data <= 8'hFF;
            16'd29402: data <= 8'h1F;
            16'd29403: data <= 8'h00;
            16'd29404: data <= 8'h1F;
            16'd29405: data <= 8'h00;
            16'd29406: data <= 8'h1F;
            16'd29407: data <= 8'h00;
            16'd29408: data <= 8'h1F;
            16'd29409: data <= 8'h00;
            16'd29410: data <= 8'h1F;
            16'd29411: data <= 8'h00;
            16'd29412: data <= 8'h1F;
            16'd29413: data <= 8'h00;
            16'd29414: data <= 8'h1F;
            16'd29415: data <= 8'h00;
            16'd29416: data <= 8'h1F;
            16'd29417: data <= 8'h00;
            16'd29418: data <= 8'h1F;
            16'd29419: data <= 8'h00;
            16'd29420: data <= 8'h1F;
            16'd29421: data <= 8'h00;
            16'd29422: data <= 8'h1F;
            16'd29423: data <= 8'h00;
            16'd29424: data <= 8'h1F;
            16'd29425: data <= 8'h00;
            16'd29426: data <= 8'h1F;
            16'd29427: data <= 8'h00;
            16'd29428: data <= 8'h1F;
            16'd29429: data <= 8'h00;
            16'd29430: data <= 8'h1F;
            16'd29431: data <= 8'h00;
            16'd29432: data <= 8'h1F;
            16'd29433: data <= 8'h00;
            16'd29434: data <= 8'h1F;
            16'd29435: data <= 8'h00;
            16'd29436: data <= 8'h1F;
            16'd29437: data <= 8'h00;
            16'd29438: data <= 8'h1F;
            16'd29439: data <= 8'h00;
            16'd29440: data <= 8'hFF;
            16'd29441: data <= 8'hFF;
            16'd29442: data <= 8'h1F;
            16'd29443: data <= 8'h00;
            16'd29444: data <= 8'h1F;
            16'd29445: data <= 8'h00;
            16'd29446: data <= 8'h1F;
            16'd29447: data <= 8'h00;
            16'd29448: data <= 8'h1F;
            16'd29449: data <= 8'h00;
            16'd29450: data <= 8'h1F;
            16'd29451: data <= 8'h00;
            16'd29452: data <= 8'h1F;
            16'd29453: data <= 8'h00;
            16'd29454: data <= 8'h1F;
            16'd29455: data <= 8'h00;
            16'd29456: data <= 8'h1F;
            16'd29457: data <= 8'h00;
            16'd29458: data <= 8'h1F;
            16'd29459: data <= 8'h00;
            16'd29460: data <= 8'h1F;
            16'd29461: data <= 8'h00;
            16'd29462: data <= 8'h1F;
            16'd29463: data <= 8'h00;
            16'd29464: data <= 8'h1F;
            16'd29465: data <= 8'h00;
            16'd29466: data <= 8'h1F;
            16'd29467: data <= 8'h00;
            16'd29468: data <= 8'h1F;
            16'd29469: data <= 8'h00;
            16'd29470: data <= 8'h1F;
            16'd29471: data <= 8'h00;
            16'd29472: data <= 8'h1F;
            16'd29473: data <= 8'h00;
            16'd29474: data <= 8'h1F;
            16'd29475: data <= 8'h00;
            16'd29476: data <= 8'h1F;
            16'd29477: data <= 8'h00;
            16'd29478: data <= 8'h1F;
            16'd29479: data <= 8'h00;
            16'd29480: data <= 8'hFF;
            16'd29481: data <= 8'hFF;
            16'd29482: data <= 8'h1F;
            16'd29483: data <= 8'h00;
            16'd29484: data <= 8'h1F;
            16'd29485: data <= 8'h00;
            16'd29486: data <= 8'h1F;
            16'd29487: data <= 8'h00;
            16'd29488: data <= 8'h1F;
            16'd29489: data <= 8'h00;
            16'd29490: data <= 8'h1F;
            16'd29491: data <= 8'h00;
            16'd29492: data <= 8'h1F;
            16'd29493: data <= 8'h00;
            16'd29494: data <= 8'h1F;
            16'd29495: data <= 8'h00;
            16'd29496: data <= 8'h1F;
            16'd29497: data <= 8'h00;
            16'd29498: data <= 8'h1F;
            16'd29499: data <= 8'h00;
            16'd29500: data <= 8'h1F;
            16'd29501: data <= 8'h00;
            16'd29502: data <= 8'h1F;
            16'd29503: data <= 8'h00;
            16'd29504: data <= 8'h1F;
            16'd29505: data <= 8'h00;
            16'd29506: data <= 8'h1F;
            16'd29507: data <= 8'h00;
            16'd29508: data <= 8'h1F;
            16'd29509: data <= 8'h00;
            16'd29510: data <= 8'h1F;
            16'd29511: data <= 8'h00;
            16'd29512: data <= 8'h1F;
            16'd29513: data <= 8'h00;
            16'd29514: data <= 8'h1F;
            16'd29515: data <= 8'h00;
            16'd29516: data <= 8'h1F;
            16'd29517: data <= 8'h00;
            16'd29518: data <= 8'h1F;
            16'd29519: data <= 8'h00;
            16'd29520: data <= 8'hFF;
            16'd29521: data <= 8'hFF;
            16'd29522: data <= 8'h1F;
            16'd29523: data <= 8'h00;
            16'd29524: data <= 8'h1F;
            16'd29525: data <= 8'h00;
            16'd29526: data <= 8'h1F;
            16'd29527: data <= 8'h00;
            16'd29528: data <= 8'h1F;
            16'd29529: data <= 8'h00;
            16'd29530: data <= 8'h1F;
            16'd29531: data <= 8'h00;
            16'd29532: data <= 8'h1F;
            16'd29533: data <= 8'h00;
            16'd29534: data <= 8'h1F;
            16'd29535: data <= 8'h00;
            16'd29536: data <= 8'h1F;
            16'd29537: data <= 8'h00;
            16'd29538: data <= 8'h1F;
            16'd29539: data <= 8'h00;
            16'd29540: data <= 8'h1F;
            16'd29541: data <= 8'h00;
            16'd29542: data <= 8'h1F;
            16'd29543: data <= 8'h00;
            16'd29544: data <= 8'h1F;
            16'd29545: data <= 8'h00;
            16'd29546: data <= 8'h1F;
            16'd29547: data <= 8'h00;
            16'd29548: data <= 8'h1F;
            16'd29549: data <= 8'h00;
            16'd29550: data <= 8'h1F;
            16'd29551: data <= 8'h00;
            16'd29552: data <= 8'h1F;
            16'd29553: data <= 8'h00;
            16'd29554: data <= 8'h1F;
            16'd29555: data <= 8'h00;
            16'd29556: data <= 8'h1F;
            16'd29557: data <= 8'h00;
            16'd29558: data <= 8'h1F;
            16'd29559: data <= 8'h00;
            16'd29560: data <= 8'hFF;
            16'd29561: data <= 8'hFF;
            16'd29562: data <= 8'h1F;
            16'd29563: data <= 8'h00;
            16'd29564: data <= 8'h1F;
            16'd29565: data <= 8'h00;
            16'd29566: data <= 8'h1F;
            16'd29567: data <= 8'h00;
            16'd29568: data <= 8'h1F;
            16'd29569: data <= 8'h00;
            16'd29570: data <= 8'h1F;
            16'd29571: data <= 8'h00;
            16'd29572: data <= 8'h1F;
            16'd29573: data <= 8'h00;
            16'd29574: data <= 8'h1F;
            16'd29575: data <= 8'h00;
            16'd29576: data <= 8'h1F;
            16'd29577: data <= 8'h00;
            16'd29578: data <= 8'h1F;
            16'd29579: data <= 8'h00;
            16'd29580: data <= 8'h1F;
            16'd29581: data <= 8'h00;
            16'd29582: data <= 8'h1F;
            16'd29583: data <= 8'h00;
            16'd29584: data <= 8'h1F;
            16'd29585: data <= 8'h00;
            16'd29586: data <= 8'h1F;
            16'd29587: data <= 8'h00;
            16'd29588: data <= 8'h1F;
            16'd29589: data <= 8'h00;
            16'd29590: data <= 8'h1F;
            16'd29591: data <= 8'h00;
            16'd29592: data <= 8'h1F;
            16'd29593: data <= 8'h00;
            16'd29594: data <= 8'h1F;
            16'd29595: data <= 8'h00;
            16'd29596: data <= 8'h1F;
            16'd29597: data <= 8'h00;
            16'd29598: data <= 8'h1F;
            16'd29599: data <= 8'h00;
            16'd29600: data <= 8'hFF;
            16'd29601: data <= 8'hFF;
            16'd29602: data <= 8'h1F;
            16'd29603: data <= 8'h00;
            16'd29604: data <= 8'h1F;
            16'd29605: data <= 8'h00;
            16'd29606: data <= 8'h1F;
            16'd29607: data <= 8'h00;
            16'd29608: data <= 8'h1F;
            16'd29609: data <= 8'h00;
            16'd29610: data <= 8'h1F;
            16'd29611: data <= 8'h00;
            16'd29612: data <= 8'h1F;
            16'd29613: data <= 8'h00;
            16'd29614: data <= 8'h1F;
            16'd29615: data <= 8'h00;
            16'd29616: data <= 8'h1F;
            16'd29617: data <= 8'h00;
            16'd29618: data <= 8'h1F;
            16'd29619: data <= 8'h00;
            16'd29620: data <= 8'h1F;
            16'd29621: data <= 8'h00;
            16'd29622: data <= 8'h1F;
            16'd29623: data <= 8'h00;
            16'd29624: data <= 8'h1F;
            16'd29625: data <= 8'h00;
            16'd29626: data <= 8'h1F;
            16'd29627: data <= 8'h00;
            16'd29628: data <= 8'h1F;
            16'd29629: data <= 8'h00;
            16'd29630: data <= 8'h1F;
            16'd29631: data <= 8'h00;
            16'd29632: data <= 8'h1F;
            16'd29633: data <= 8'h00;
            16'd29634: data <= 8'h1F;
            16'd29635: data <= 8'h00;
            16'd29636: data <= 8'h1F;
            16'd29637: data <= 8'h00;
            16'd29638: data <= 8'h1F;
            16'd29639: data <= 8'h00;
            16'd29640: data <= 8'hFF;
            16'd29641: data <= 8'hFF;
            16'd29642: data <= 8'h1F;
            16'd29643: data <= 8'h00;
            16'd29644: data <= 8'h1F;
            16'd29645: data <= 8'h00;
            16'd29646: data <= 8'h1F;
            16'd29647: data <= 8'h00;
            16'd29648: data <= 8'h1F;
            16'd29649: data <= 8'h00;
            16'd29650: data <= 8'h1F;
            16'd29651: data <= 8'h00;
            16'd29652: data <= 8'h1F;
            16'd29653: data <= 8'h00;
            16'd29654: data <= 8'h1F;
            16'd29655: data <= 8'h00;
            16'd29656: data <= 8'h1F;
            16'd29657: data <= 8'h00;
            16'd29658: data <= 8'h1F;
            16'd29659: data <= 8'h00;
            16'd29660: data <= 8'h1F;
            16'd29661: data <= 8'h00;
            16'd29662: data <= 8'h1F;
            16'd29663: data <= 8'h00;
            16'd29664: data <= 8'h1F;
            16'd29665: data <= 8'h00;
            16'd29666: data <= 8'h1F;
            16'd29667: data <= 8'h00;
            16'd29668: data <= 8'h1F;
            16'd29669: data <= 8'h00;
            16'd29670: data <= 8'h1F;
            16'd29671: data <= 8'h00;
            16'd29672: data <= 8'h1F;
            16'd29673: data <= 8'h00;
            16'd29674: data <= 8'h1F;
            16'd29675: data <= 8'h00;
            16'd29676: data <= 8'h1F;
            16'd29677: data <= 8'h00;
            16'd29678: data <= 8'h1F;
            16'd29679: data <= 8'h00;
            16'd29680: data <= 8'hFF;
            16'd29681: data <= 8'hFF;
            16'd29682: data <= 8'h1F;
            16'd29683: data <= 8'h00;
            16'd29684: data <= 8'h1F;
            16'd29685: data <= 8'h00;
            16'd29686: data <= 8'h1F;
            16'd29687: data <= 8'h00;
            16'd29688: data <= 8'h1F;
            16'd29689: data <= 8'h00;
            16'd29690: data <= 8'h1F;
            16'd29691: data <= 8'h00;
            16'd29692: data <= 8'h1F;
            16'd29693: data <= 8'h00;
            16'd29694: data <= 8'h1F;
            16'd29695: data <= 8'h00;
            16'd29696: data <= 8'h1F;
            16'd29697: data <= 8'h00;
            16'd29698: data <= 8'h1F;
            16'd29699: data <= 8'h00;
            16'd29700: data <= 8'h1F;
            16'd29701: data <= 8'h00;
            16'd29702: data <= 8'h1F;
            16'd29703: data <= 8'h00;
            16'd29704: data <= 8'h1F;
            16'd29705: data <= 8'h00;
            16'd29706: data <= 8'h1F;
            16'd29707: data <= 8'h00;
            16'd29708: data <= 8'h1F;
            16'd29709: data <= 8'h00;
            16'd29710: data <= 8'h1F;
            16'd29711: data <= 8'h00;
            16'd29712: data <= 8'h1F;
            16'd29713: data <= 8'h00;
            16'd29714: data <= 8'h1F;
            16'd29715: data <= 8'h00;
            16'd29716: data <= 8'h1F;
            16'd29717: data <= 8'h00;
            16'd29718: data <= 8'h1F;
            16'd29719: data <= 8'h00;
            16'd29720: data <= 8'hFF;
            16'd29721: data <= 8'hFF;
            16'd29722: data <= 8'h1F;
            16'd29723: data <= 8'h00;
            16'd29724: data <= 8'h1F;
            16'd29725: data <= 8'h00;
            16'd29726: data <= 8'h1F;
            16'd29727: data <= 8'h00;
            16'd29728: data <= 8'h1F;
            16'd29729: data <= 8'h00;
            16'd29730: data <= 8'h1F;
            16'd29731: data <= 8'h00;
            16'd29732: data <= 8'h1F;
            16'd29733: data <= 8'h00;
            16'd29734: data <= 8'h1F;
            16'd29735: data <= 8'h00;
            16'd29736: data <= 8'h1F;
            16'd29737: data <= 8'h00;
            16'd29738: data <= 8'h1F;
            16'd29739: data <= 8'h00;
            16'd29740: data <= 8'h1F;
            16'd29741: data <= 8'h00;
            16'd29742: data <= 8'h1F;
            16'd29743: data <= 8'h00;
            16'd29744: data <= 8'h1F;
            16'd29745: data <= 8'h00;
            16'd29746: data <= 8'h1F;
            16'd29747: data <= 8'h00;
            16'd29748: data <= 8'h1F;
            16'd29749: data <= 8'h00;
            16'd29750: data <= 8'h1F;
            16'd29751: data <= 8'h00;
            16'd29752: data <= 8'h1F;
            16'd29753: data <= 8'h00;
            16'd29754: data <= 8'h1F;
            16'd29755: data <= 8'h00;
            16'd29756: data <= 8'h1F;
            16'd29757: data <= 8'h00;
            16'd29758: data <= 8'h1F;
            16'd29759: data <= 8'h00;
            16'd29760: data <= 8'hFF;
            16'd29761: data <= 8'hFF;
            16'd29762: data <= 8'h1F;
            16'd29763: data <= 8'h00;
            16'd29764: data <= 8'h1F;
            16'd29765: data <= 8'h00;
            16'd29766: data <= 8'h1F;
            16'd29767: data <= 8'h00;
            16'd29768: data <= 8'h1F;
            16'd29769: data <= 8'h00;
            16'd29770: data <= 8'h1F;
            16'd29771: data <= 8'h00;
            16'd29772: data <= 8'h1F;
            16'd29773: data <= 8'h00;
            16'd29774: data <= 8'h1F;
            16'd29775: data <= 8'h00;
            16'd29776: data <= 8'h1F;
            16'd29777: data <= 8'h00;
            16'd29778: data <= 8'h1F;
            16'd29779: data <= 8'h00;
            16'd29780: data <= 8'h1F;
            16'd29781: data <= 8'h00;
            16'd29782: data <= 8'h1F;
            16'd29783: data <= 8'h00;
            16'd29784: data <= 8'h1F;
            16'd29785: data <= 8'h00;
            16'd29786: data <= 8'h1F;
            16'd29787: data <= 8'h00;
            16'd29788: data <= 8'h1F;
            16'd29789: data <= 8'h00;
            16'd29790: data <= 8'h1F;
            16'd29791: data <= 8'h00;
            16'd29792: data <= 8'h1F;
            16'd29793: data <= 8'h00;
            16'd29794: data <= 8'h1F;
            16'd29795: data <= 8'h00;
            16'd29796: data <= 8'h1F;
            16'd29797: data <= 8'h00;
            16'd29798: data <= 8'h1F;
            16'd29799: data <= 8'h00;
            16'd29800: data <= 8'hFF;
            16'd29801: data <= 8'hFF;
            16'd29802: data <= 8'h1F;
            16'd29803: data <= 8'h00;
            16'd29804: data <= 8'h1F;
            16'd29805: data <= 8'h00;
            16'd29806: data <= 8'h1F;
            16'd29807: data <= 8'h00;
            16'd29808: data <= 8'h1F;
            16'd29809: data <= 8'h00;
            16'd29810: data <= 8'h1F;
            16'd29811: data <= 8'h00;
            16'd29812: data <= 8'h1F;
            16'd29813: data <= 8'h00;
            16'd29814: data <= 8'h1F;
            16'd29815: data <= 8'h00;
            16'd29816: data <= 8'h1F;
            16'd29817: data <= 8'h00;
            16'd29818: data <= 8'h1F;
            16'd29819: data <= 8'h00;
            16'd29820: data <= 8'h1F;
            16'd29821: data <= 8'h00;
            16'd29822: data <= 8'h1F;
            16'd29823: data <= 8'h00;
            16'd29824: data <= 8'h1F;
            16'd29825: data <= 8'h00;
            16'd29826: data <= 8'h1F;
            16'd29827: data <= 8'h00;
            16'd29828: data <= 8'h1F;
            16'd29829: data <= 8'h00;
            16'd29830: data <= 8'h1F;
            16'd29831: data <= 8'h00;
            16'd29832: data <= 8'h1F;
            16'd29833: data <= 8'h00;
            16'd29834: data <= 8'h1F;
            16'd29835: data <= 8'h00;
            16'd29836: data <= 8'h1F;
            16'd29837: data <= 8'h00;
            16'd29838: data <= 8'h1F;
            16'd29839: data <= 8'h00;
            16'd29840: data <= 8'hFF;
            16'd29841: data <= 8'hFF;
            16'd29842: data <= 8'h1F;
            16'd29843: data <= 8'h00;
            16'd29844: data <= 8'h1F;
            16'd29845: data <= 8'h00;
            16'd29846: data <= 8'h1F;
            16'd29847: data <= 8'h00;
            16'd29848: data <= 8'h1F;
            16'd29849: data <= 8'h00;
            16'd29850: data <= 8'h1F;
            16'd29851: data <= 8'h00;
            16'd29852: data <= 8'h1F;
            16'd29853: data <= 8'h00;
            16'd29854: data <= 8'h1F;
            16'd29855: data <= 8'h00;
            16'd29856: data <= 8'h1F;
            16'd29857: data <= 8'h00;
            16'd29858: data <= 8'h1F;
            16'd29859: data <= 8'h00;
            16'd29860: data <= 8'h1F;
            16'd29861: data <= 8'h00;
            16'd29862: data <= 8'h1F;
            16'd29863: data <= 8'h00;
            16'd29864: data <= 8'h1F;
            16'd29865: data <= 8'h00;
            16'd29866: data <= 8'h1F;
            16'd29867: data <= 8'h00;
            16'd29868: data <= 8'h1F;
            16'd29869: data <= 8'h00;
            16'd29870: data <= 8'h1F;
            16'd29871: data <= 8'h00;
            16'd29872: data <= 8'h1F;
            16'd29873: data <= 8'h00;
            16'd29874: data <= 8'h1F;
            16'd29875: data <= 8'h00;
            16'd29876: data <= 8'h1F;
            16'd29877: data <= 8'h00;
            16'd29878: data <= 8'h1F;
            16'd29879: data <= 8'h00;
            16'd29880: data <= 8'hFF;
            16'd29881: data <= 8'hFF;
            16'd29882: data <= 8'h1F;
            16'd29883: data <= 8'h00;
            16'd29884: data <= 8'h1F;
            16'd29885: data <= 8'h00;
            16'd29886: data <= 8'h1F;
            16'd29887: data <= 8'h00;
            16'd29888: data <= 8'h1F;
            16'd29889: data <= 8'h00;
            16'd29890: data <= 8'h1F;
            16'd29891: data <= 8'h00;
            16'd29892: data <= 8'h1F;
            16'd29893: data <= 8'h00;
            16'd29894: data <= 8'h1F;
            16'd29895: data <= 8'h00;
            16'd29896: data <= 8'h1F;
            16'd29897: data <= 8'h00;
            16'd29898: data <= 8'h1F;
            16'd29899: data <= 8'h00;
            16'd29900: data <= 8'h1F;
            16'd29901: data <= 8'h00;
            16'd29902: data <= 8'h1F;
            16'd29903: data <= 8'h00;
            16'd29904: data <= 8'h1F;
            16'd29905: data <= 8'h00;
            16'd29906: data <= 8'h1F;
            16'd29907: data <= 8'h00;
            16'd29908: data <= 8'h1F;
            16'd29909: data <= 8'h00;
            16'd29910: data <= 8'h1F;
            16'd29911: data <= 8'h00;
            16'd29912: data <= 8'h1F;
            16'd29913: data <= 8'h00;
            16'd29914: data <= 8'h1F;
            16'd29915: data <= 8'h00;
            16'd29916: data <= 8'h1F;
            16'd29917: data <= 8'h00;
            16'd29918: data <= 8'h1F;
            16'd29919: data <= 8'h00;
            16'd29920: data <= 8'hFF;
            16'd29921: data <= 8'hFF;
            16'd29922: data <= 8'h1F;
            16'd29923: data <= 8'h00;
            16'd29924: data <= 8'h1F;
            16'd29925: data <= 8'h00;
            16'd29926: data <= 8'h1F;
            16'd29927: data <= 8'h00;
            16'd29928: data <= 8'h1F;
            16'd29929: data <= 8'h00;
            16'd29930: data <= 8'h1F;
            16'd29931: data <= 8'h00;
            16'd29932: data <= 8'h1F;
            16'd29933: data <= 8'h00;
            16'd29934: data <= 8'h1F;
            16'd29935: data <= 8'h00;
            16'd29936: data <= 8'h1F;
            16'd29937: data <= 8'h00;
            16'd29938: data <= 8'h1F;
            16'd29939: data <= 8'h00;
            16'd29940: data <= 8'h1F;
            16'd29941: data <= 8'h00;
            16'd29942: data <= 8'h1F;
            16'd29943: data <= 8'h00;
            16'd29944: data <= 8'h1F;
            16'd29945: data <= 8'h00;
            16'd29946: data <= 8'h1F;
            16'd29947: data <= 8'h00;
            16'd29948: data <= 8'h1F;
            16'd29949: data <= 8'h00;
            16'd29950: data <= 8'h1F;
            16'd29951: data <= 8'h00;
            16'd29952: data <= 8'h1F;
            16'd29953: data <= 8'h00;
            16'd29954: data <= 8'h1F;
            16'd29955: data <= 8'h00;
            16'd29956: data <= 8'h1F;
            16'd29957: data <= 8'h00;
            16'd29958: data <= 8'h1F;
            16'd29959: data <= 8'h00;
            16'd29960: data <= 8'hFF;
            16'd29961: data <= 8'hFF;
            16'd29962: data <= 8'h1F;
            16'd29963: data <= 8'h00;
            16'd29964: data <= 8'h1F;
            16'd29965: data <= 8'h00;
            16'd29966: data <= 8'h1F;
            16'd29967: data <= 8'h00;
            16'd29968: data <= 8'h1F;
            16'd29969: data <= 8'h00;
            16'd29970: data <= 8'h1F;
            16'd29971: data <= 8'h00;
            16'd29972: data <= 8'h1F;
            16'd29973: data <= 8'h00;
            16'd29974: data <= 8'h1F;
            16'd29975: data <= 8'h00;
            16'd29976: data <= 8'h1F;
            16'd29977: data <= 8'h00;
            16'd29978: data <= 8'h1F;
            16'd29979: data <= 8'h00;
            16'd29980: data <= 8'h1F;
            16'd29981: data <= 8'h00;
            16'd29982: data <= 8'h1F;
            16'd29983: data <= 8'h00;
            16'd29984: data <= 8'h1F;
            16'd29985: data <= 8'h00;
            16'd29986: data <= 8'h1F;
            16'd29987: data <= 8'h00;
            16'd29988: data <= 8'h1F;
            16'd29989: data <= 8'h00;
            16'd29990: data <= 8'h1F;
            16'd29991: data <= 8'h00;
            16'd29992: data <= 8'h1F;
            16'd29993: data <= 8'h00;
            16'd29994: data <= 8'h1F;
            16'd29995: data <= 8'h00;
            16'd29996: data <= 8'h1F;
            16'd29997: data <= 8'h00;
            16'd29998: data <= 8'h1F;
            16'd29999: data <= 8'h00;
            16'd30000: data <= 8'hFF;
            16'd30001: data <= 8'hFF;
            16'd30002: data <= 8'h1F;
            16'd30003: data <= 8'h00;
            16'd30004: data <= 8'h1F;
            16'd30005: data <= 8'h00;
            16'd30006: data <= 8'h1F;
            16'd30007: data <= 8'h00;
            16'd30008: data <= 8'h1F;
            16'd30009: data <= 8'h00;
            16'd30010: data <= 8'h1F;
            16'd30011: data <= 8'h00;
            16'd30012: data <= 8'h1F;
            16'd30013: data <= 8'h00;
            16'd30014: data <= 8'h1F;
            16'd30015: data <= 8'h00;
            16'd30016: data <= 8'h1F;
            16'd30017: data <= 8'h00;
            16'd30018: data <= 8'h1F;
            16'd30019: data <= 8'h00;
            16'd30020: data <= 8'h1F;
            16'd30021: data <= 8'h00;
            16'd30022: data <= 8'h1F;
            16'd30023: data <= 8'h00;
            16'd30024: data <= 8'h1F;
            16'd30025: data <= 8'h00;
            16'd30026: data <= 8'h1F;
            16'd30027: data <= 8'h00;
            16'd30028: data <= 8'h1F;
            16'd30029: data <= 8'h00;
            16'd30030: data <= 8'h1F;
            16'd30031: data <= 8'h00;
            16'd30032: data <= 8'h1F;
            16'd30033: data <= 8'h00;
            16'd30034: data <= 8'h1F;
            16'd30035: data <= 8'h00;
            16'd30036: data <= 8'h1F;
            16'd30037: data <= 8'h00;
            16'd30038: data <= 8'h1F;
            16'd30039: data <= 8'h00;
            16'd30040: data <= 8'hFF;
            16'd30041: data <= 8'hFF;
            16'd30042: data <= 8'h1F;
            16'd30043: data <= 8'h00;
            16'd30044: data <= 8'h1F;
            16'd30045: data <= 8'h00;
            16'd30046: data <= 8'h1F;
            16'd30047: data <= 8'h00;
            16'd30048: data <= 8'h1F;
            16'd30049: data <= 8'h00;
            16'd30050: data <= 8'h1F;
            16'd30051: data <= 8'h00;
            16'd30052: data <= 8'h1F;
            16'd30053: data <= 8'h00;
            16'd30054: data <= 8'h1F;
            16'd30055: data <= 8'h00;
            16'd30056: data <= 8'h1F;
            16'd30057: data <= 8'h00;
            16'd30058: data <= 8'h1F;
            16'd30059: data <= 8'h00;
            16'd30060: data <= 8'h1F;
            16'd30061: data <= 8'h00;
            16'd30062: data <= 8'h1F;
            16'd30063: data <= 8'h00;
            16'd30064: data <= 8'h1F;
            16'd30065: data <= 8'h00;
            16'd30066: data <= 8'h1F;
            16'd30067: data <= 8'h00;
            16'd30068: data <= 8'h1F;
            16'd30069: data <= 8'h00;
            16'd30070: data <= 8'h1F;
            16'd30071: data <= 8'h00;
            16'd30072: data <= 8'h1F;
            16'd30073: data <= 8'h00;
            16'd30074: data <= 8'h1F;
            16'd30075: data <= 8'h00;
            16'd30076: data <= 8'h1F;
            16'd30077: data <= 8'h00;
            16'd30078: data <= 8'h1F;
            16'd30079: data <= 8'h00;
            16'd30080: data <= 8'hFF;
            16'd30081: data <= 8'hFF;
            16'd30082: data <= 8'h1F;
            16'd30083: data <= 8'h00;
            16'd30084: data <= 8'h1F;
            16'd30085: data <= 8'h00;
            16'd30086: data <= 8'h1F;
            16'd30087: data <= 8'h00;
            16'd30088: data <= 8'h1F;
            16'd30089: data <= 8'h00;
            16'd30090: data <= 8'h1F;
            16'd30091: data <= 8'h00;
            16'd30092: data <= 8'h1F;
            16'd30093: data <= 8'h00;
            16'd30094: data <= 8'h1F;
            16'd30095: data <= 8'h00;
            16'd30096: data <= 8'h1F;
            16'd30097: data <= 8'h00;
            16'd30098: data <= 8'h1F;
            16'd30099: data <= 8'h00;
            16'd30100: data <= 8'h1F;
            16'd30101: data <= 8'h00;
            16'd30102: data <= 8'h1F;
            16'd30103: data <= 8'h00;
            16'd30104: data <= 8'h1F;
            16'd30105: data <= 8'h00;
            16'd30106: data <= 8'h1F;
            16'd30107: data <= 8'h00;
            16'd30108: data <= 8'h1F;
            16'd30109: data <= 8'h00;
            16'd30110: data <= 8'h1F;
            16'd30111: data <= 8'h00;
            16'd30112: data <= 8'h1F;
            16'd30113: data <= 8'h00;
            16'd30114: data <= 8'h1F;
            16'd30115: data <= 8'h00;
            16'd30116: data <= 8'h1F;
            16'd30117: data <= 8'h00;
            16'd30118: data <= 8'h1F;
            16'd30119: data <= 8'h00;
            16'd30120: data <= 8'hFF;
            16'd30121: data <= 8'hFF;
            16'd30122: data <= 8'h1F;
            16'd30123: data <= 8'h00;
            16'd30124: data <= 8'h1F;
            16'd30125: data <= 8'h00;
            16'd30126: data <= 8'h1F;
            16'd30127: data <= 8'h00;
            16'd30128: data <= 8'h1F;
            16'd30129: data <= 8'h00;
            16'd30130: data <= 8'h1F;
            16'd30131: data <= 8'h00;
            16'd30132: data <= 8'h1F;
            16'd30133: data <= 8'h00;
            16'd30134: data <= 8'h1F;
            16'd30135: data <= 8'h00;
            16'd30136: data <= 8'h1F;
            16'd30137: data <= 8'h00;
            16'd30138: data <= 8'h1F;
            16'd30139: data <= 8'h00;
            16'd30140: data <= 8'h1F;
            16'd30141: data <= 8'h00;
            16'd30142: data <= 8'h1F;
            16'd30143: data <= 8'h00;
            16'd30144: data <= 8'h1F;
            16'd30145: data <= 8'h00;
            16'd30146: data <= 8'h1F;
            16'd30147: data <= 8'h00;
            16'd30148: data <= 8'h1F;
            16'd30149: data <= 8'h00;
            16'd30150: data <= 8'h1F;
            16'd30151: data <= 8'h00;
            16'd30152: data <= 8'h1F;
            16'd30153: data <= 8'h00;
            16'd30154: data <= 8'h1F;
            16'd30155: data <= 8'h00;
            16'd30156: data <= 8'h1F;
            16'd30157: data <= 8'h00;
            16'd30158: data <= 8'h1F;
            16'd30159: data <= 8'h00;
            16'd30160: data <= 8'hFF;
            16'd30161: data <= 8'hFF;
            16'd30162: data <= 8'h1F;
            16'd30163: data <= 8'h00;
            16'd30164: data <= 8'h1F;
            16'd30165: data <= 8'h00;
            16'd30166: data <= 8'h1F;
            16'd30167: data <= 8'h00;
            16'd30168: data <= 8'h1F;
            16'd30169: data <= 8'h00;
            16'd30170: data <= 8'h1F;
            16'd30171: data <= 8'h00;
            16'd30172: data <= 8'h1F;
            16'd30173: data <= 8'h00;
            16'd30174: data <= 8'h1F;
            16'd30175: data <= 8'h00;
            16'd30176: data <= 8'h1F;
            16'd30177: data <= 8'h00;
            16'd30178: data <= 8'h1F;
            16'd30179: data <= 8'h00;
            16'd30180: data <= 8'h1F;
            16'd30181: data <= 8'h00;
            16'd30182: data <= 8'h1F;
            16'd30183: data <= 8'h00;
            16'd30184: data <= 8'h1F;
            16'd30185: data <= 8'h00;
            16'd30186: data <= 8'h1F;
            16'd30187: data <= 8'h00;
            16'd30188: data <= 8'h1F;
            16'd30189: data <= 8'h00;
            16'd30190: data <= 8'h1F;
            16'd30191: data <= 8'h00;
            16'd30192: data <= 8'h1F;
            16'd30193: data <= 8'h00;
            16'd30194: data <= 8'h1F;
            16'd30195: data <= 8'h00;
            16'd30196: data <= 8'h1F;
            16'd30197: data <= 8'h00;
            16'd30198: data <= 8'h1F;
            16'd30199: data <= 8'h00;
            16'd30200: data <= 8'hFF;
            16'd30201: data <= 8'hFF;
            16'd30202: data <= 8'h1F;
            16'd30203: data <= 8'h00;
            16'd30204: data <= 8'h1F;
            16'd30205: data <= 8'h00;
            16'd30206: data <= 8'h1F;
            16'd30207: data <= 8'h00;
            16'd30208: data <= 8'h1F;
            16'd30209: data <= 8'h00;
            16'd30210: data <= 8'h1F;
            16'd30211: data <= 8'h00;
            16'd30212: data <= 8'h1F;
            16'd30213: data <= 8'h00;
            16'd30214: data <= 8'h1F;
            16'd30215: data <= 8'h00;
            16'd30216: data <= 8'h1F;
            16'd30217: data <= 8'h00;
            16'd30218: data <= 8'h1F;
            16'd30219: data <= 8'h00;
            16'd30220: data <= 8'h1F;
            16'd30221: data <= 8'h00;
            16'd30222: data <= 8'h1F;
            16'd30223: data <= 8'h00;
            16'd30224: data <= 8'h1F;
            16'd30225: data <= 8'h00;
            16'd30226: data <= 8'h1F;
            16'd30227: data <= 8'h00;
            16'd30228: data <= 8'h1F;
            16'd30229: data <= 8'h00;
            16'd30230: data <= 8'h1F;
            16'd30231: data <= 8'h00;
            16'd30232: data <= 8'h1F;
            16'd30233: data <= 8'h00;
            16'd30234: data <= 8'h1F;
            16'd30235: data <= 8'h00;
            16'd30236: data <= 8'h1F;
            16'd30237: data <= 8'h00;
            16'd30238: data <= 8'h1F;
            16'd30239: data <= 8'h00;
            16'd30240: data <= 8'hFF;
            16'd30241: data <= 8'hFF;
            16'd30242: data <= 8'h1F;
            16'd30243: data <= 8'h00;
            16'd30244: data <= 8'h1F;
            16'd30245: data <= 8'h00;
            16'd30246: data <= 8'h1F;
            16'd30247: data <= 8'h00;
            16'd30248: data <= 8'h1F;
            16'd30249: data <= 8'h00;
            16'd30250: data <= 8'h1F;
            16'd30251: data <= 8'h00;
            16'd30252: data <= 8'h1F;
            16'd30253: data <= 8'h00;
            16'd30254: data <= 8'h1F;
            16'd30255: data <= 8'h00;
            16'd30256: data <= 8'h1F;
            16'd30257: data <= 8'h00;
            16'd30258: data <= 8'h1F;
            16'd30259: data <= 8'h00;
            16'd30260: data <= 8'h1F;
            16'd30261: data <= 8'h00;
            16'd30262: data <= 8'h1F;
            16'd30263: data <= 8'h00;
            16'd30264: data <= 8'h1F;
            16'd30265: data <= 8'h00;
            16'd30266: data <= 8'h1F;
            16'd30267: data <= 8'h00;
            16'd30268: data <= 8'h1F;
            16'd30269: data <= 8'h00;
            16'd30270: data <= 8'h1F;
            16'd30271: data <= 8'h00;
            16'd30272: data <= 8'h1F;
            16'd30273: data <= 8'h00;
            16'd30274: data <= 8'h1F;
            16'd30275: data <= 8'h00;
            16'd30276: data <= 8'h1F;
            16'd30277: data <= 8'h00;
            16'd30278: data <= 8'h1F;
            16'd30279: data <= 8'h00;
            16'd30280: data <= 8'hFF;
            16'd30281: data <= 8'hFF;
            16'd30282: data <= 8'h1F;
            16'd30283: data <= 8'h00;
            16'd30284: data <= 8'h1F;
            16'd30285: data <= 8'h00;
            16'd30286: data <= 8'h1F;
            16'd30287: data <= 8'h00;
            16'd30288: data <= 8'h1F;
            16'd30289: data <= 8'h00;
            16'd30290: data <= 8'h1F;
            16'd30291: data <= 8'h00;
            16'd30292: data <= 8'h1F;
            16'd30293: data <= 8'h00;
            16'd30294: data <= 8'h1F;
            16'd30295: data <= 8'h00;
            16'd30296: data <= 8'h1F;
            16'd30297: data <= 8'h00;
            16'd30298: data <= 8'h1F;
            16'd30299: data <= 8'h00;
            16'd30300: data <= 8'h1F;
            16'd30301: data <= 8'h00;
            16'd30302: data <= 8'h1F;
            16'd30303: data <= 8'h00;
            16'd30304: data <= 8'h1F;
            16'd30305: data <= 8'h00;
            16'd30306: data <= 8'h1F;
            16'd30307: data <= 8'h00;
            16'd30308: data <= 8'h1F;
            16'd30309: data <= 8'h00;
            16'd30310: data <= 8'h1F;
            16'd30311: data <= 8'h00;
            16'd30312: data <= 8'h1F;
            16'd30313: data <= 8'h00;
            16'd30314: data <= 8'h1F;
            16'd30315: data <= 8'h00;
            16'd30316: data <= 8'h1F;
            16'd30317: data <= 8'h00;
            16'd30318: data <= 8'h1F;
            16'd30319: data <= 8'h00;
            16'd30320: data <= 8'hFF;
            16'd30321: data <= 8'hFF;
            16'd30322: data <= 8'h1F;
            16'd30323: data <= 8'h00;
            16'd30324: data <= 8'h1F;
            16'd30325: data <= 8'h00;
            16'd30326: data <= 8'h1F;
            16'd30327: data <= 8'h00;
            16'd30328: data <= 8'h1F;
            16'd30329: data <= 8'h00;
            16'd30330: data <= 8'h1F;
            16'd30331: data <= 8'h00;
            16'd30332: data <= 8'h1F;
            16'd30333: data <= 8'h00;
            16'd30334: data <= 8'h1F;
            16'd30335: data <= 8'h00;
            16'd30336: data <= 8'h1F;
            16'd30337: data <= 8'h00;
            16'd30338: data <= 8'h1F;
            16'd30339: data <= 8'h00;
            16'd30340: data <= 8'h1F;
            16'd30341: data <= 8'h00;
            16'd30342: data <= 8'h1F;
            16'd30343: data <= 8'h00;
            16'd30344: data <= 8'h1F;
            16'd30345: data <= 8'h00;
            16'd30346: data <= 8'h1F;
            16'd30347: data <= 8'h00;
            16'd30348: data <= 8'h1F;
            16'd30349: data <= 8'h00;
            16'd30350: data <= 8'h1F;
            16'd30351: data <= 8'h00;
            16'd30352: data <= 8'h1F;
            16'd30353: data <= 8'h00;
            16'd30354: data <= 8'h1F;
            16'd30355: data <= 8'h00;
            16'd30356: data <= 8'h1F;
            16'd30357: data <= 8'h00;
            16'd30358: data <= 8'h1F;
            16'd30359: data <= 8'h00;
            16'd30360: data <= 8'hFF;
            16'd30361: data <= 8'hFF;
            16'd30362: data <= 8'h1F;
            16'd30363: data <= 8'h00;
            16'd30364: data <= 8'h1F;
            16'd30365: data <= 8'h00;
            16'd30366: data <= 8'h1F;
            16'd30367: data <= 8'h00;
            16'd30368: data <= 8'h1F;
            16'd30369: data <= 8'h00;
            16'd30370: data <= 8'h1F;
            16'd30371: data <= 8'h00;
            16'd30372: data <= 8'h1F;
            16'd30373: data <= 8'h00;
            16'd30374: data <= 8'h1F;
            16'd30375: data <= 8'h00;
            16'd30376: data <= 8'h1F;
            16'd30377: data <= 8'h00;
            16'd30378: data <= 8'h1F;
            16'd30379: data <= 8'h00;
            16'd30380: data <= 8'h1F;
            16'd30381: data <= 8'h00;
            16'd30382: data <= 8'h1F;
            16'd30383: data <= 8'h00;
            16'd30384: data <= 8'h1F;
            16'd30385: data <= 8'h00;
            16'd30386: data <= 8'h1F;
            16'd30387: data <= 8'h00;
            16'd30388: data <= 8'h1F;
            16'd30389: data <= 8'h00;
            16'd30390: data <= 8'h1F;
            16'd30391: data <= 8'h00;
            16'd30392: data <= 8'h1F;
            16'd30393: data <= 8'h00;
            16'd30394: data <= 8'h1F;
            16'd30395: data <= 8'h00;
            16'd30396: data <= 8'h1F;
            16'd30397: data <= 8'h00;
            16'd30398: data <= 8'h1F;
            16'd30399: data <= 8'h00;
            16'd30400: data <= 8'hFF;
            16'd30401: data <= 8'hFF;
            16'd30402: data <= 8'h1F;
            16'd30403: data <= 8'h00;
            16'd30404: data <= 8'h1F;
            16'd30405: data <= 8'h00;
            16'd30406: data <= 8'h1F;
            16'd30407: data <= 8'h00;
            16'd30408: data <= 8'h1F;
            16'd30409: data <= 8'h00;
            16'd30410: data <= 8'h1F;
            16'd30411: data <= 8'h00;
            16'd30412: data <= 8'h1F;
            16'd30413: data <= 8'h00;
            16'd30414: data <= 8'h1F;
            16'd30415: data <= 8'h00;
            16'd30416: data <= 8'h1F;
            16'd30417: data <= 8'h00;
            16'd30418: data <= 8'h1F;
            16'd30419: data <= 8'h00;
            16'd30420: data <= 8'h1F;
            16'd30421: data <= 8'h00;
            16'd30422: data <= 8'h1F;
            16'd30423: data <= 8'h00;
            16'd30424: data <= 8'h1F;
            16'd30425: data <= 8'h00;
            16'd30426: data <= 8'h1F;
            16'd30427: data <= 8'h00;
            16'd30428: data <= 8'h1F;
            16'd30429: data <= 8'h00;
            16'd30430: data <= 8'h1F;
            16'd30431: data <= 8'h00;
            16'd30432: data <= 8'h1F;
            16'd30433: data <= 8'h00;
            16'd30434: data <= 8'h1F;
            16'd30435: data <= 8'h00;
            16'd30436: data <= 8'h1F;
            16'd30437: data <= 8'h00;
            16'd30438: data <= 8'h1F;
            16'd30439: data <= 8'h00;
            16'd30440: data <= 8'hFF;
            16'd30441: data <= 8'hFF;
            16'd30442: data <= 8'h1F;
            16'd30443: data <= 8'h00;
            16'd30444: data <= 8'h1F;
            16'd30445: data <= 8'h00;
            16'd30446: data <= 8'h1F;
            16'd30447: data <= 8'h00;
            16'd30448: data <= 8'h1F;
            16'd30449: data <= 8'h00;
            16'd30450: data <= 8'h1F;
            16'd30451: data <= 8'h00;
            16'd30452: data <= 8'h1F;
            16'd30453: data <= 8'h00;
            16'd30454: data <= 8'h1F;
            16'd30455: data <= 8'h00;
            16'd30456: data <= 8'h1F;
            16'd30457: data <= 8'h00;
            16'd30458: data <= 8'h1F;
            16'd30459: data <= 8'h00;
            16'd30460: data <= 8'h1F;
            16'd30461: data <= 8'h00;
            16'd30462: data <= 8'h1F;
            16'd30463: data <= 8'h00;
            16'd30464: data <= 8'h1F;
            16'd30465: data <= 8'h00;
            16'd30466: data <= 8'h1F;
            16'd30467: data <= 8'h00;
            16'd30468: data <= 8'h1F;
            16'd30469: data <= 8'h00;
            16'd30470: data <= 8'h1F;
            16'd30471: data <= 8'h00;
            16'd30472: data <= 8'h1F;
            16'd30473: data <= 8'h00;
            16'd30474: data <= 8'h1F;
            16'd30475: data <= 8'h00;
            16'd30476: data <= 8'h1F;
            16'd30477: data <= 8'h00;
            16'd30478: data <= 8'h1F;
            16'd30479: data <= 8'h00;
            16'd30480: data <= 8'hFF;
            16'd30481: data <= 8'hFF;
            16'd30482: data <= 8'h1F;
            16'd30483: data <= 8'h00;
            16'd30484: data <= 8'h1F;
            16'd30485: data <= 8'h00;
            16'd30486: data <= 8'h1F;
            16'd30487: data <= 8'h00;
            16'd30488: data <= 8'h1F;
            16'd30489: data <= 8'h00;
            16'd30490: data <= 8'h1F;
            16'd30491: data <= 8'h00;
            16'd30492: data <= 8'h1F;
            16'd30493: data <= 8'h00;
            16'd30494: data <= 8'h1F;
            16'd30495: data <= 8'h00;
            16'd30496: data <= 8'h1F;
            16'd30497: data <= 8'h00;
            16'd30498: data <= 8'h1F;
            16'd30499: data <= 8'h00;
            16'd30500: data <= 8'h1F;
            16'd30501: data <= 8'h00;
            16'd30502: data <= 8'h1F;
            16'd30503: data <= 8'h00;
            16'd30504: data <= 8'h1F;
            16'd30505: data <= 8'h00;
            16'd30506: data <= 8'h1F;
            16'd30507: data <= 8'h00;
            16'd30508: data <= 8'h1F;
            16'd30509: data <= 8'h00;
            16'd30510: data <= 8'h1F;
            16'd30511: data <= 8'h00;
            16'd30512: data <= 8'h1F;
            16'd30513: data <= 8'h00;
            16'd30514: data <= 8'h1F;
            16'd30515: data <= 8'h00;
            16'd30516: data <= 8'h1F;
            16'd30517: data <= 8'h00;
            16'd30518: data <= 8'h1F;
            16'd30519: data <= 8'h00;
            16'd30520: data <= 8'hFF;
            16'd30521: data <= 8'hFF;
            16'd30522: data <= 8'h1F;
            16'd30523: data <= 8'h00;
            16'd30524: data <= 8'h1F;
            16'd30525: data <= 8'h00;
            16'd30526: data <= 8'h1F;
            16'd30527: data <= 8'h00;
            16'd30528: data <= 8'h1F;
            16'd30529: data <= 8'h00;
            16'd30530: data <= 8'h1F;
            16'd30531: data <= 8'h00;
            16'd30532: data <= 8'h1F;
            16'd30533: data <= 8'h00;
            16'd30534: data <= 8'h1F;
            16'd30535: data <= 8'h00;
            16'd30536: data <= 8'h1F;
            16'd30537: data <= 8'h00;
            16'd30538: data <= 8'h1F;
            16'd30539: data <= 8'h00;
            16'd30540: data <= 8'h1F;
            16'd30541: data <= 8'h00;
            16'd30542: data <= 8'h1F;
            16'd30543: data <= 8'h00;
            16'd30544: data <= 8'h1F;
            16'd30545: data <= 8'h00;
            16'd30546: data <= 8'h1F;
            16'd30547: data <= 8'h00;
            16'd30548: data <= 8'h1F;
            16'd30549: data <= 8'h00;
            16'd30550: data <= 8'h1F;
            16'd30551: data <= 8'h00;
            16'd30552: data <= 8'h1F;
            16'd30553: data <= 8'h00;
            16'd30554: data <= 8'h1F;
            16'd30555: data <= 8'h00;
            16'd30556: data <= 8'h1F;
            16'd30557: data <= 8'h00;
            16'd30558: data <= 8'h1F;
            16'd30559: data <= 8'h00;
            16'd30560: data <= 8'hFF;
            16'd30561: data <= 8'hFF;
            16'd30562: data <= 8'h1F;
            16'd30563: data <= 8'h00;
            16'd30564: data <= 8'h1F;
            16'd30565: data <= 8'h00;
            16'd30566: data <= 8'h1F;
            16'd30567: data <= 8'h00;
            16'd30568: data <= 8'h1F;
            16'd30569: data <= 8'h00;
            16'd30570: data <= 8'h1F;
            16'd30571: data <= 8'h00;
            16'd30572: data <= 8'h1F;
            16'd30573: data <= 8'h00;
            16'd30574: data <= 8'h1F;
            16'd30575: data <= 8'h00;
            16'd30576: data <= 8'h1F;
            16'd30577: data <= 8'h00;
            16'd30578: data <= 8'h1F;
            16'd30579: data <= 8'h00;
            16'd30580: data <= 8'h1F;
            16'd30581: data <= 8'h00;
            16'd30582: data <= 8'h1F;
            16'd30583: data <= 8'h00;
            16'd30584: data <= 8'h1F;
            16'd30585: data <= 8'h00;
            16'd30586: data <= 8'h1F;
            16'd30587: data <= 8'h00;
            16'd30588: data <= 8'h1F;
            16'd30589: data <= 8'h00;
            16'd30590: data <= 8'h1F;
            16'd30591: data <= 8'h00;
            16'd30592: data <= 8'h1F;
            16'd30593: data <= 8'h00;
            16'd30594: data <= 8'h1F;
            16'd30595: data <= 8'h00;
            16'd30596: data <= 8'h1F;
            16'd30597: data <= 8'h00;
            16'd30598: data <= 8'h1F;
            16'd30599: data <= 8'h00;
            16'd30600: data <= 8'hFF;
            16'd30601: data <= 8'hFF;
            16'd30602: data <= 8'h1F;
            16'd30603: data <= 8'h00;
            16'd30604: data <= 8'h1F;
            16'd30605: data <= 8'h00;
            16'd30606: data <= 8'h1F;
            16'd30607: data <= 8'h00;
            16'd30608: data <= 8'h1F;
            16'd30609: data <= 8'h00;
            16'd30610: data <= 8'h1F;
            16'd30611: data <= 8'h00;
            16'd30612: data <= 8'h1F;
            16'd30613: data <= 8'h00;
            16'd30614: data <= 8'h1F;
            16'd30615: data <= 8'h00;
            16'd30616: data <= 8'h1F;
            16'd30617: data <= 8'h00;
            16'd30618: data <= 8'h1F;
            16'd30619: data <= 8'h00;
            16'd30620: data <= 8'h1F;
            16'd30621: data <= 8'h00;
            16'd30622: data <= 8'h1F;
            16'd30623: data <= 8'h00;
            16'd30624: data <= 8'h1F;
            16'd30625: data <= 8'h00;
            16'd30626: data <= 8'h1F;
            16'd30627: data <= 8'h00;
            16'd30628: data <= 8'h1F;
            16'd30629: data <= 8'h00;
            16'd30630: data <= 8'h1F;
            16'd30631: data <= 8'h00;
            16'd30632: data <= 8'h1F;
            16'd30633: data <= 8'h00;
            16'd30634: data <= 8'h1F;
            16'd30635: data <= 8'h00;
            16'd30636: data <= 8'h1F;
            16'd30637: data <= 8'h00;
            16'd30638: data <= 8'h1F;
            16'd30639: data <= 8'h00;
            16'd30640: data <= 8'hFF;
            16'd30641: data <= 8'hFF;
            16'd30642: data <= 8'h1F;
            16'd30643: data <= 8'h00;
            16'd30644: data <= 8'h1F;
            16'd30645: data <= 8'h00;
            16'd30646: data <= 8'h1F;
            16'd30647: data <= 8'h00;
            16'd30648: data <= 8'h1F;
            16'd30649: data <= 8'h00;
            16'd30650: data <= 8'h1F;
            16'd30651: data <= 8'h00;
            16'd30652: data <= 8'h1F;
            16'd30653: data <= 8'h00;
            16'd30654: data <= 8'h1F;
            16'd30655: data <= 8'h00;
            16'd30656: data <= 8'h1F;
            16'd30657: data <= 8'h00;
            16'd30658: data <= 8'h1F;
            16'd30659: data <= 8'h00;
            16'd30660: data <= 8'h1F;
            16'd30661: data <= 8'h00;
            16'd30662: data <= 8'h1F;
            16'd30663: data <= 8'h00;
            16'd30664: data <= 8'h1F;
            16'd30665: data <= 8'h00;
            16'd30666: data <= 8'h1F;
            16'd30667: data <= 8'h00;
            16'd30668: data <= 8'h1F;
            16'd30669: data <= 8'h00;
            16'd30670: data <= 8'h1F;
            16'd30671: data <= 8'h00;
            16'd30672: data <= 8'h1F;
            16'd30673: data <= 8'h00;
            16'd30674: data <= 8'h1F;
            16'd30675: data <= 8'h00;
            16'd30676: data <= 8'h1F;
            16'd30677: data <= 8'h00;
            16'd30678: data <= 8'h1F;
            16'd30679: data <= 8'h00;
            16'd30680: data <= 8'hFF;
            16'd30681: data <= 8'hFF;
            16'd30682: data <= 8'h1F;
            16'd30683: data <= 8'h00;
            16'd30684: data <= 8'h1F;
            16'd30685: data <= 8'h00;
            16'd30686: data <= 8'h1F;
            16'd30687: data <= 8'h00;
            16'd30688: data <= 8'h1F;
            16'd30689: data <= 8'h00;
            16'd30690: data <= 8'h1F;
            16'd30691: data <= 8'h00;
            16'd30692: data <= 8'h1F;
            16'd30693: data <= 8'h00;
            16'd30694: data <= 8'h1F;
            16'd30695: data <= 8'h00;
            16'd30696: data <= 8'h1F;
            16'd30697: data <= 8'h00;
            16'd30698: data <= 8'h1F;
            16'd30699: data <= 8'h00;
            16'd30700: data <= 8'h1F;
            16'd30701: data <= 8'h00;
            16'd30702: data <= 8'h1F;
            16'd30703: data <= 8'h00;
            16'd30704: data <= 8'h1F;
            16'd30705: data <= 8'h00;
            16'd30706: data <= 8'h1F;
            16'd30707: data <= 8'h00;
            16'd30708: data <= 8'h1F;
            16'd30709: data <= 8'h00;
            16'd30710: data <= 8'h1F;
            16'd30711: data <= 8'h00;
            16'd30712: data <= 8'h1F;
            16'd30713: data <= 8'h00;
            16'd30714: data <= 8'h1F;
            16'd30715: data <= 8'h00;
            16'd30716: data <= 8'h1F;
            16'd30717: data <= 8'h00;
            16'd30718: data <= 8'h1F;
            16'd30719: data <= 8'h00;
            16'd30720: data <= 8'hFF;
            16'd30721: data <= 8'hFF;
            16'd30722: data <= 8'h1F;
            16'd30723: data <= 8'h00;
            16'd30724: data <= 8'h1F;
            16'd30725: data <= 8'h00;
            16'd30726: data <= 8'h1F;
            16'd30727: data <= 8'h00;
            16'd30728: data <= 8'h1F;
            16'd30729: data <= 8'h00;
            16'd30730: data <= 8'h1F;
            16'd30731: data <= 8'h00;
            16'd30732: data <= 8'h1F;
            16'd30733: data <= 8'h00;
            16'd30734: data <= 8'h1F;
            16'd30735: data <= 8'h00;
            16'd30736: data <= 8'h1F;
            16'd30737: data <= 8'h00;
            16'd30738: data <= 8'h1F;
            16'd30739: data <= 8'h00;
            16'd30740: data <= 8'h1F;
            16'd30741: data <= 8'h00;
            16'd30742: data <= 8'h1F;
            16'd30743: data <= 8'h00;
            16'd30744: data <= 8'h1F;
            16'd30745: data <= 8'h00;
            16'd30746: data <= 8'h1F;
            16'd30747: data <= 8'h00;
            16'd30748: data <= 8'h1F;
            16'd30749: data <= 8'h00;
            16'd30750: data <= 8'h1F;
            16'd30751: data <= 8'h00;
            16'd30752: data <= 8'h1F;
            16'd30753: data <= 8'h00;
            16'd30754: data <= 8'h1F;
            16'd30755: data <= 8'h00;
            16'd30756: data <= 8'h1F;
            16'd30757: data <= 8'h00;
            16'd30758: data <= 8'h1F;
            16'd30759: data <= 8'h00;
            16'd30760: data <= 8'hFF;
            16'd30761: data <= 8'hFF;
            16'd30762: data <= 8'h1F;
            16'd30763: data <= 8'h00;
            16'd30764: data <= 8'h1F;
            16'd30765: data <= 8'h00;
            16'd30766: data <= 8'h1F;
            16'd30767: data <= 8'h00;
            16'd30768: data <= 8'h1F;
            16'd30769: data <= 8'h00;
            16'd30770: data <= 8'h1F;
            16'd30771: data <= 8'h00;
            16'd30772: data <= 8'h1F;
            16'd30773: data <= 8'h00;
            16'd30774: data <= 8'h1F;
            16'd30775: data <= 8'h00;
            16'd30776: data <= 8'h1F;
            16'd30777: data <= 8'h00;
            16'd30778: data <= 8'h1F;
            16'd30779: data <= 8'h00;
            16'd30780: data <= 8'h1F;
            16'd30781: data <= 8'h00;
            16'd30782: data <= 8'h1F;
            16'd30783: data <= 8'h00;
            16'd30784: data <= 8'h1F;
            16'd30785: data <= 8'h00;
            16'd30786: data <= 8'h1F;
            16'd30787: data <= 8'h00;
            16'd30788: data <= 8'h1F;
            16'd30789: data <= 8'h00;
            16'd30790: data <= 8'h1F;
            16'd30791: data <= 8'h00;
            16'd30792: data <= 8'h1F;
            16'd30793: data <= 8'h00;
            16'd30794: data <= 8'h1F;
            16'd30795: data <= 8'h00;
            16'd30796: data <= 8'h1F;
            16'd30797: data <= 8'h00;
            16'd30798: data <= 8'h1F;
            16'd30799: data <= 8'h00;
            16'd30800: data <= 8'hFF;
            16'd30801: data <= 8'hFF;
            16'd30802: data <= 8'h1F;
            16'd30803: data <= 8'h00;
            16'd30804: data <= 8'h1F;
            16'd30805: data <= 8'h00;
            16'd30806: data <= 8'h1F;
            16'd30807: data <= 8'h00;
            16'd30808: data <= 8'h1F;
            16'd30809: data <= 8'h00;
            16'd30810: data <= 8'h1F;
            16'd30811: data <= 8'h00;
            16'd30812: data <= 8'h1F;
            16'd30813: data <= 8'h00;
            16'd30814: data <= 8'h1F;
            16'd30815: data <= 8'h00;
            16'd30816: data <= 8'h1F;
            16'd30817: data <= 8'h00;
            16'd30818: data <= 8'h1F;
            16'd30819: data <= 8'h00;
            16'd30820: data <= 8'h1F;
            16'd30821: data <= 8'h00;
            16'd30822: data <= 8'h1F;
            16'd30823: data <= 8'h00;
            16'd30824: data <= 8'h1F;
            16'd30825: data <= 8'h00;
            16'd30826: data <= 8'h1F;
            16'd30827: data <= 8'h00;
            16'd30828: data <= 8'h1F;
            16'd30829: data <= 8'h00;
            16'd30830: data <= 8'h1F;
            16'd30831: data <= 8'h00;
            16'd30832: data <= 8'h1F;
            16'd30833: data <= 8'h00;
            16'd30834: data <= 8'h1F;
            16'd30835: data <= 8'h00;
            16'd30836: data <= 8'h1F;
            16'd30837: data <= 8'h00;
            16'd30838: data <= 8'h1F;
            16'd30839: data <= 8'h00;
            16'd30840: data <= 8'hFF;
            16'd30841: data <= 8'hFF;
            16'd30842: data <= 8'h1F;
            16'd30843: data <= 8'h00;
            16'd30844: data <= 8'h1F;
            16'd30845: data <= 8'h00;
            16'd30846: data <= 8'h1F;
            16'd30847: data <= 8'h00;
            16'd30848: data <= 8'h1F;
            16'd30849: data <= 8'h00;
            16'd30850: data <= 8'h1F;
            16'd30851: data <= 8'h00;
            16'd30852: data <= 8'h1F;
            16'd30853: data <= 8'h00;
            16'd30854: data <= 8'h1F;
            16'd30855: data <= 8'h00;
            16'd30856: data <= 8'h1F;
            16'd30857: data <= 8'h00;
            16'd30858: data <= 8'h1F;
            16'd30859: data <= 8'h00;
            16'd30860: data <= 8'h1F;
            16'd30861: data <= 8'h00;
            16'd30862: data <= 8'h1F;
            16'd30863: data <= 8'h00;
            16'd30864: data <= 8'h1F;
            16'd30865: data <= 8'h00;
            16'd30866: data <= 8'h1F;
            16'd30867: data <= 8'h00;
            16'd30868: data <= 8'h1F;
            16'd30869: data <= 8'h00;
            16'd30870: data <= 8'h1F;
            16'd30871: data <= 8'h00;
            16'd30872: data <= 8'h1F;
            16'd30873: data <= 8'h00;
            16'd30874: data <= 8'h1F;
            16'd30875: data <= 8'h00;
            16'd30876: data <= 8'h1F;
            16'd30877: data <= 8'h00;
            16'd30878: data <= 8'h1F;
            16'd30879: data <= 8'h00;
            16'd30880: data <= 8'hFF;
            16'd30881: data <= 8'hFF;
            16'd30882: data <= 8'h1F;
            16'd30883: data <= 8'h00;
            16'd30884: data <= 8'h1F;
            16'd30885: data <= 8'h00;
            16'd30886: data <= 8'h1F;
            16'd30887: data <= 8'h00;
            16'd30888: data <= 8'h1F;
            16'd30889: data <= 8'h00;
            16'd30890: data <= 8'h1F;
            16'd30891: data <= 8'h00;
            16'd30892: data <= 8'h1F;
            16'd30893: data <= 8'h00;
            16'd30894: data <= 8'h1F;
            16'd30895: data <= 8'h00;
            16'd30896: data <= 8'h1F;
            16'd30897: data <= 8'h00;
            16'd30898: data <= 8'h1F;
            16'd30899: data <= 8'h00;
            16'd30900: data <= 8'h1F;
            16'd30901: data <= 8'h00;
            16'd30902: data <= 8'h1F;
            16'd30903: data <= 8'h00;
            16'd30904: data <= 8'h1F;
            16'd30905: data <= 8'h00;
            16'd30906: data <= 8'h1F;
            16'd30907: data <= 8'h00;
            16'd30908: data <= 8'h1F;
            16'd30909: data <= 8'h00;
            16'd30910: data <= 8'h1F;
            16'd30911: data <= 8'h00;
            16'd30912: data <= 8'h1F;
            16'd30913: data <= 8'h00;
            16'd30914: data <= 8'h1F;
            16'd30915: data <= 8'h00;
            16'd30916: data <= 8'h1F;
            16'd30917: data <= 8'h00;
            16'd30918: data <= 8'h1F;
            16'd30919: data <= 8'h00;
            16'd30920: data <= 8'hFF;
            16'd30921: data <= 8'hFF;
            16'd30922: data <= 8'h1F;
            16'd30923: data <= 8'h00;
            16'd30924: data <= 8'h1F;
            16'd30925: data <= 8'h00;
            16'd30926: data <= 8'h1F;
            16'd30927: data <= 8'h00;
            16'd30928: data <= 8'h1F;
            16'd30929: data <= 8'h00;
            16'd30930: data <= 8'h1F;
            16'd30931: data <= 8'h00;
            16'd30932: data <= 8'h1F;
            16'd30933: data <= 8'h00;
            16'd30934: data <= 8'h1F;
            16'd30935: data <= 8'h00;
            16'd30936: data <= 8'h1F;
            16'd30937: data <= 8'h00;
            16'd30938: data <= 8'h1F;
            16'd30939: data <= 8'h00;
            16'd30940: data <= 8'h1F;
            16'd30941: data <= 8'h00;
            16'd30942: data <= 8'h1F;
            16'd30943: data <= 8'h00;
            16'd30944: data <= 8'h1F;
            16'd30945: data <= 8'h00;
            16'd30946: data <= 8'h1F;
            16'd30947: data <= 8'h00;
            16'd30948: data <= 8'h1F;
            16'd30949: data <= 8'h00;
            16'd30950: data <= 8'h1F;
            16'd30951: data <= 8'h00;
            16'd30952: data <= 8'h1F;
            16'd30953: data <= 8'h00;
            16'd30954: data <= 8'h1F;
            16'd30955: data <= 8'h00;
            16'd30956: data <= 8'h1F;
            16'd30957: data <= 8'h00;
            16'd30958: data <= 8'h1F;
            16'd30959: data <= 8'h00;
            16'd30960: data <= 8'hFF;
            16'd30961: data <= 8'hFF;
            16'd30962: data <= 8'h1F;
            16'd30963: data <= 8'h00;
            16'd30964: data <= 8'h1F;
            16'd30965: data <= 8'h00;
            16'd30966: data <= 8'h1F;
            16'd30967: data <= 8'h00;
            16'd30968: data <= 8'h1F;
            16'd30969: data <= 8'h00;
            16'd30970: data <= 8'h1F;
            16'd30971: data <= 8'h00;
            16'd30972: data <= 8'h1F;
            16'd30973: data <= 8'h00;
            16'd30974: data <= 8'h1F;
            16'd30975: data <= 8'h00;
            16'd30976: data <= 8'h1F;
            16'd30977: data <= 8'h00;
            16'd30978: data <= 8'h1F;
            16'd30979: data <= 8'h00;
            16'd30980: data <= 8'h1F;
            16'd30981: data <= 8'h00;
            16'd30982: data <= 8'h1F;
            16'd30983: data <= 8'h00;
            16'd30984: data <= 8'h1F;
            16'd30985: data <= 8'h00;
            16'd30986: data <= 8'h1F;
            16'd30987: data <= 8'h00;
            16'd30988: data <= 8'h1F;
            16'd30989: data <= 8'h00;
            16'd30990: data <= 8'h1F;
            16'd30991: data <= 8'h00;
            16'd30992: data <= 8'h1F;
            16'd30993: data <= 8'h00;
            16'd30994: data <= 8'h1F;
            16'd30995: data <= 8'h00;
            16'd30996: data <= 8'h1F;
            16'd30997: data <= 8'h00;
            16'd30998: data <= 8'h1F;
            16'd30999: data <= 8'h00;
            16'd31000: data <= 8'hFF;
            16'd31001: data <= 8'hFF;
            16'd31002: data <= 8'h1F;
            16'd31003: data <= 8'h00;
            16'd31004: data <= 8'h1F;
            16'd31005: data <= 8'h00;
            16'd31006: data <= 8'h1F;
            16'd31007: data <= 8'h00;
            16'd31008: data <= 8'h1F;
            16'd31009: data <= 8'h00;
            16'd31010: data <= 8'h1F;
            16'd31011: data <= 8'h00;
            16'd31012: data <= 8'h1F;
            16'd31013: data <= 8'h00;
            16'd31014: data <= 8'h1F;
            16'd31015: data <= 8'h00;
            16'd31016: data <= 8'h1F;
            16'd31017: data <= 8'h00;
            16'd31018: data <= 8'h1F;
            16'd31019: data <= 8'h00;
            16'd31020: data <= 8'h1F;
            16'd31021: data <= 8'h00;
            16'd31022: data <= 8'h1F;
            16'd31023: data <= 8'h00;
            16'd31024: data <= 8'h1F;
            16'd31025: data <= 8'h00;
            16'd31026: data <= 8'h1F;
            16'd31027: data <= 8'h00;
            16'd31028: data <= 8'h1F;
            16'd31029: data <= 8'h00;
            16'd31030: data <= 8'h1F;
            16'd31031: data <= 8'h00;
            16'd31032: data <= 8'h1F;
            16'd31033: data <= 8'h00;
            16'd31034: data <= 8'h1F;
            16'd31035: data <= 8'h00;
            16'd31036: data <= 8'h1F;
            16'd31037: data <= 8'h00;
            16'd31038: data <= 8'h1F;
            16'd31039: data <= 8'h00;
            16'd31040: data <= 8'hFF;
            16'd31041: data <= 8'hFF;
            16'd31042: data <= 8'h1F;
            16'd31043: data <= 8'h00;
            16'd31044: data <= 8'h1F;
            16'd31045: data <= 8'h00;
            16'd31046: data <= 8'h1F;
            16'd31047: data <= 8'h00;
            16'd31048: data <= 8'h1F;
            16'd31049: data <= 8'h00;
            16'd31050: data <= 8'h1F;
            16'd31051: data <= 8'h00;
            16'd31052: data <= 8'h1F;
            16'd31053: data <= 8'h00;
            16'd31054: data <= 8'h1F;
            16'd31055: data <= 8'h00;
            16'd31056: data <= 8'h1F;
            16'd31057: data <= 8'h00;
            16'd31058: data <= 8'h1F;
            16'd31059: data <= 8'h00;
            16'd31060: data <= 8'h1F;
            16'd31061: data <= 8'h00;
            16'd31062: data <= 8'h1F;
            16'd31063: data <= 8'h00;
            16'd31064: data <= 8'h1F;
            16'd31065: data <= 8'h00;
            16'd31066: data <= 8'h1F;
            16'd31067: data <= 8'h00;
            16'd31068: data <= 8'h1F;
            16'd31069: data <= 8'h00;
            16'd31070: data <= 8'h1F;
            16'd31071: data <= 8'h00;
            16'd31072: data <= 8'h1F;
            16'd31073: data <= 8'h00;
            16'd31074: data <= 8'h1F;
            16'd31075: data <= 8'h00;
            16'd31076: data <= 8'h1F;
            16'd31077: data <= 8'h00;
            16'd31078: data <= 8'h1F;
            16'd31079: data <= 8'h00;
            16'd31080: data <= 8'hFF;
            16'd31081: data <= 8'hFF;
            16'd31082: data <= 8'h1F;
            16'd31083: data <= 8'h00;
            16'd31084: data <= 8'h1F;
            16'd31085: data <= 8'h00;
            16'd31086: data <= 8'h1F;
            16'd31087: data <= 8'h00;
            16'd31088: data <= 8'h1F;
            16'd31089: data <= 8'h00;
            16'd31090: data <= 8'h1F;
            16'd31091: data <= 8'h00;
            16'd31092: data <= 8'h1F;
            16'd31093: data <= 8'h00;
            16'd31094: data <= 8'h1F;
            16'd31095: data <= 8'h00;
            16'd31096: data <= 8'h1F;
            16'd31097: data <= 8'h00;
            16'd31098: data <= 8'h1F;
            16'd31099: data <= 8'h00;
            16'd31100: data <= 8'h1F;
            16'd31101: data <= 8'h00;
            16'd31102: data <= 8'h1F;
            16'd31103: data <= 8'h00;
            16'd31104: data <= 8'h1F;
            16'd31105: data <= 8'h00;
            16'd31106: data <= 8'h1F;
            16'd31107: data <= 8'h00;
            16'd31108: data <= 8'h1F;
            16'd31109: data <= 8'h00;
            16'd31110: data <= 8'h1F;
            16'd31111: data <= 8'h00;
            16'd31112: data <= 8'h1F;
            16'd31113: data <= 8'h00;
            16'd31114: data <= 8'h1F;
            16'd31115: data <= 8'h00;
            16'd31116: data <= 8'h1F;
            16'd31117: data <= 8'h00;
            16'd31118: data <= 8'h1F;
            16'd31119: data <= 8'h00;
            16'd31120: data <= 8'hFF;
            16'd31121: data <= 8'hFF;
            16'd31122: data <= 8'h1F;
            16'd31123: data <= 8'h00;
            16'd31124: data <= 8'h1F;
            16'd31125: data <= 8'h00;
            16'd31126: data <= 8'h1F;
            16'd31127: data <= 8'h00;
            16'd31128: data <= 8'h1F;
            16'd31129: data <= 8'h00;
            16'd31130: data <= 8'h1F;
            16'd31131: data <= 8'h00;
            16'd31132: data <= 8'h1F;
            16'd31133: data <= 8'h00;
            16'd31134: data <= 8'h1F;
            16'd31135: data <= 8'h00;
            16'd31136: data <= 8'h1F;
            16'd31137: data <= 8'h00;
            16'd31138: data <= 8'h1F;
            16'd31139: data <= 8'h00;
            16'd31140: data <= 8'h1F;
            16'd31141: data <= 8'h00;
            16'd31142: data <= 8'h1F;
            16'd31143: data <= 8'h00;
            16'd31144: data <= 8'h1F;
            16'd31145: data <= 8'h00;
            16'd31146: data <= 8'h1F;
            16'd31147: data <= 8'h00;
            16'd31148: data <= 8'h1F;
            16'd31149: data <= 8'h00;
            16'd31150: data <= 8'h1F;
            16'd31151: data <= 8'h00;
            16'd31152: data <= 8'h1F;
            16'd31153: data <= 8'h00;
            16'd31154: data <= 8'h1F;
            16'd31155: data <= 8'h00;
            16'd31156: data <= 8'h1F;
            16'd31157: data <= 8'h00;
            16'd31158: data <= 8'h1F;
            16'd31159: data <= 8'h00;
            16'd31160: data <= 8'hFF;
            16'd31161: data <= 8'hFF;
            16'd31162: data <= 8'h1F;
            16'd31163: data <= 8'h00;
            16'd31164: data <= 8'h1F;
            16'd31165: data <= 8'h00;
            16'd31166: data <= 8'h1F;
            16'd31167: data <= 8'h00;
            16'd31168: data <= 8'h1F;
            16'd31169: data <= 8'h00;
            16'd31170: data <= 8'h1F;
            16'd31171: data <= 8'h00;
            16'd31172: data <= 8'h1F;
            16'd31173: data <= 8'h00;
            16'd31174: data <= 8'h1F;
            16'd31175: data <= 8'h00;
            16'd31176: data <= 8'h1F;
            16'd31177: data <= 8'h00;
            16'd31178: data <= 8'h1F;
            16'd31179: data <= 8'h00;
            16'd31180: data <= 8'h1F;
            16'd31181: data <= 8'h00;
            16'd31182: data <= 8'h1F;
            16'd31183: data <= 8'h00;
            16'd31184: data <= 8'h1F;
            16'd31185: data <= 8'h00;
            16'd31186: data <= 8'h1F;
            16'd31187: data <= 8'h00;
            16'd31188: data <= 8'h1F;
            16'd31189: data <= 8'h00;
            16'd31190: data <= 8'h1F;
            16'd31191: data <= 8'h00;
            16'd31192: data <= 8'h1F;
            16'd31193: data <= 8'h00;
            16'd31194: data <= 8'h1F;
            16'd31195: data <= 8'h00;
            16'd31196: data <= 8'h1F;
            16'd31197: data <= 8'h00;
            16'd31198: data <= 8'h1F;
            16'd31199: data <= 8'h00;
            16'd31200: data <= 8'hFF;
            16'd31201: data <= 8'hFF;
            16'd31202: data <= 8'h1F;
            16'd31203: data <= 8'h00;
            16'd31204: data <= 8'h1F;
            16'd31205: data <= 8'h00;
            16'd31206: data <= 8'h1F;
            16'd31207: data <= 8'h00;
            16'd31208: data <= 8'h1F;
            16'd31209: data <= 8'h00;
            16'd31210: data <= 8'h1F;
            16'd31211: data <= 8'h00;
            16'd31212: data <= 8'h1F;
            16'd31213: data <= 8'h00;
            16'd31214: data <= 8'h1F;
            16'd31215: data <= 8'h00;
            16'd31216: data <= 8'h1F;
            16'd31217: data <= 8'h00;
            16'd31218: data <= 8'h1F;
            16'd31219: data <= 8'h00;
            16'd31220: data <= 8'h1F;
            16'd31221: data <= 8'h00;
            16'd31222: data <= 8'h1F;
            16'd31223: data <= 8'h00;
            16'd31224: data <= 8'h1F;
            16'd31225: data <= 8'h00;
            16'd31226: data <= 8'h1F;
            16'd31227: data <= 8'h00;
            16'd31228: data <= 8'h1F;
            16'd31229: data <= 8'h00;
            16'd31230: data <= 8'h1F;
            16'd31231: data <= 8'h00;
            16'd31232: data <= 8'h1F;
            16'd31233: data <= 8'h00;
            16'd31234: data <= 8'h1F;
            16'd31235: data <= 8'h00;
            16'd31236: data <= 8'h1F;
            16'd31237: data <= 8'h00;
            16'd31238: data <= 8'h1F;
            16'd31239: data <= 8'h00;
            16'd31240: data <= 8'hFF;
            16'd31241: data <= 8'hFF;
            16'd31242: data <= 8'h1F;
            16'd31243: data <= 8'h00;
            16'd31244: data <= 8'h1F;
            16'd31245: data <= 8'h00;
            16'd31246: data <= 8'h1F;
            16'd31247: data <= 8'h00;
            16'd31248: data <= 8'h1F;
            16'd31249: data <= 8'h00;
            16'd31250: data <= 8'h1F;
            16'd31251: data <= 8'h00;
            16'd31252: data <= 8'h1F;
            16'd31253: data <= 8'h00;
            16'd31254: data <= 8'h1F;
            16'd31255: data <= 8'h00;
            16'd31256: data <= 8'h1F;
            16'd31257: data <= 8'h00;
            16'd31258: data <= 8'h1F;
            16'd31259: data <= 8'h00;
            16'd31260: data <= 8'h1F;
            16'd31261: data <= 8'h00;
            16'd31262: data <= 8'h1F;
            16'd31263: data <= 8'h00;
            16'd31264: data <= 8'h1F;
            16'd31265: data <= 8'h00;
            16'd31266: data <= 8'h1F;
            16'd31267: data <= 8'h00;
            16'd31268: data <= 8'h1F;
            16'd31269: data <= 8'h00;
            16'd31270: data <= 8'h1F;
            16'd31271: data <= 8'h00;
            16'd31272: data <= 8'h1F;
            16'd31273: data <= 8'h00;
            16'd31274: data <= 8'h1F;
            16'd31275: data <= 8'h00;
            16'd31276: data <= 8'h1F;
            16'd31277: data <= 8'h00;
            16'd31278: data <= 8'h1F;
            16'd31279: data <= 8'h00;
            16'd31280: data <= 8'hFF;
            16'd31281: data <= 8'hFF;
            16'd31282: data <= 8'h1F;
            16'd31283: data <= 8'h00;
            16'd31284: data <= 8'h1F;
            16'd31285: data <= 8'h00;
            16'd31286: data <= 8'h1F;
            16'd31287: data <= 8'h00;
            16'd31288: data <= 8'h1F;
            16'd31289: data <= 8'h00;
            16'd31290: data <= 8'h1F;
            16'd31291: data <= 8'h00;
            16'd31292: data <= 8'h1F;
            16'd31293: data <= 8'h00;
            16'd31294: data <= 8'h1F;
            16'd31295: data <= 8'h00;
            16'd31296: data <= 8'h1F;
            16'd31297: data <= 8'h00;
            16'd31298: data <= 8'h1F;
            16'd31299: data <= 8'h00;
            16'd31300: data <= 8'h1F;
            16'd31301: data <= 8'h00;
            16'd31302: data <= 8'h1F;
            16'd31303: data <= 8'h00;
            16'd31304: data <= 8'h1F;
            16'd31305: data <= 8'h00;
            16'd31306: data <= 8'h1F;
            16'd31307: data <= 8'h00;
            16'd31308: data <= 8'h1F;
            16'd31309: data <= 8'h00;
            16'd31310: data <= 8'h1F;
            16'd31311: data <= 8'h00;
            16'd31312: data <= 8'h1F;
            16'd31313: data <= 8'h00;
            16'd31314: data <= 8'h1F;
            16'd31315: data <= 8'h00;
            16'd31316: data <= 8'h1F;
            16'd31317: data <= 8'h00;
            16'd31318: data <= 8'h1F;
            16'd31319: data <= 8'h00;
            16'd31320: data <= 8'hFF;
            16'd31321: data <= 8'hFF;
            16'd31322: data <= 8'h1F;
            16'd31323: data <= 8'h00;
            16'd31324: data <= 8'h1F;
            16'd31325: data <= 8'h00;
            16'd31326: data <= 8'h1F;
            16'd31327: data <= 8'h00;
            16'd31328: data <= 8'h1F;
            16'd31329: data <= 8'h00;
            16'd31330: data <= 8'h1F;
            16'd31331: data <= 8'h00;
            16'd31332: data <= 8'h1F;
            16'd31333: data <= 8'h00;
            16'd31334: data <= 8'h1F;
            16'd31335: data <= 8'h00;
            16'd31336: data <= 8'h1F;
            16'd31337: data <= 8'h00;
            16'd31338: data <= 8'h1F;
            16'd31339: data <= 8'h00;
            16'd31340: data <= 8'h1F;
            16'd31341: data <= 8'h00;
            16'd31342: data <= 8'h1F;
            16'd31343: data <= 8'h00;
            16'd31344: data <= 8'h1F;
            16'd31345: data <= 8'h00;
            16'd31346: data <= 8'h1F;
            16'd31347: data <= 8'h00;
            16'd31348: data <= 8'h1F;
            16'd31349: data <= 8'h00;
            16'd31350: data <= 8'h1F;
            16'd31351: data <= 8'h00;
            16'd31352: data <= 8'h1F;
            16'd31353: data <= 8'h00;
            16'd31354: data <= 8'h1F;
            16'd31355: data <= 8'h00;
            16'd31356: data <= 8'h1F;
            16'd31357: data <= 8'h00;
            16'd31358: data <= 8'h1F;
            16'd31359: data <= 8'h00;
            16'd31360: data <= 8'hFF;
            16'd31361: data <= 8'hFF;
            16'd31362: data <= 8'h1F;
            16'd31363: data <= 8'h00;
            16'd31364: data <= 8'h1F;
            16'd31365: data <= 8'h00;
            16'd31366: data <= 8'h1F;
            16'd31367: data <= 8'h00;
            16'd31368: data <= 8'h1F;
            16'd31369: data <= 8'h00;
            16'd31370: data <= 8'h1F;
            16'd31371: data <= 8'h00;
            16'd31372: data <= 8'h1F;
            16'd31373: data <= 8'h00;
            16'd31374: data <= 8'h1F;
            16'd31375: data <= 8'h00;
            16'd31376: data <= 8'h1F;
            16'd31377: data <= 8'h00;
            16'd31378: data <= 8'h1F;
            16'd31379: data <= 8'h00;
            16'd31380: data <= 8'h1F;
            16'd31381: data <= 8'h00;
            16'd31382: data <= 8'h1F;
            16'd31383: data <= 8'h00;
            16'd31384: data <= 8'h1F;
            16'd31385: data <= 8'h00;
            16'd31386: data <= 8'h1F;
            16'd31387: data <= 8'h00;
            16'd31388: data <= 8'h1F;
            16'd31389: data <= 8'h00;
            16'd31390: data <= 8'h1F;
            16'd31391: data <= 8'h00;
            16'd31392: data <= 8'h1F;
            16'd31393: data <= 8'h00;
            16'd31394: data <= 8'h1F;
            16'd31395: data <= 8'h00;
            16'd31396: data <= 8'h1F;
            16'd31397: data <= 8'h00;
            16'd31398: data <= 8'h1F;
            16'd31399: data <= 8'h00;
            16'd31400: data <= 8'hFF;
            16'd31401: data <= 8'hFF;
            16'd31402: data <= 8'h1F;
            16'd31403: data <= 8'h00;
            16'd31404: data <= 8'h1F;
            16'd31405: data <= 8'h00;
            16'd31406: data <= 8'h1F;
            16'd31407: data <= 8'h00;
            16'd31408: data <= 8'h1F;
            16'd31409: data <= 8'h00;
            16'd31410: data <= 8'h1F;
            16'd31411: data <= 8'h00;
            16'd31412: data <= 8'h1F;
            16'd31413: data <= 8'h00;
            16'd31414: data <= 8'h1F;
            16'd31415: data <= 8'h00;
            16'd31416: data <= 8'h1F;
            16'd31417: data <= 8'h00;
            16'd31418: data <= 8'h1F;
            16'd31419: data <= 8'h00;
            16'd31420: data <= 8'h1F;
            16'd31421: data <= 8'h00;
            16'd31422: data <= 8'h1F;
            16'd31423: data <= 8'h00;
            16'd31424: data <= 8'h1F;
            16'd31425: data <= 8'h00;
            16'd31426: data <= 8'h1F;
            16'd31427: data <= 8'h00;
            16'd31428: data <= 8'h1F;
            16'd31429: data <= 8'h00;
            16'd31430: data <= 8'h1F;
            16'd31431: data <= 8'h00;
            16'd31432: data <= 8'h1F;
            16'd31433: data <= 8'h00;
            16'd31434: data <= 8'h1F;
            16'd31435: data <= 8'h00;
            16'd31436: data <= 8'h1F;
            16'd31437: data <= 8'h00;
            16'd31438: data <= 8'h1F;
            16'd31439: data <= 8'h00;
            16'd31440: data <= 8'hFF;
            16'd31441: data <= 8'hFF;
            16'd31442: data <= 8'h1F;
            16'd31443: data <= 8'h00;
            16'd31444: data <= 8'h1F;
            16'd31445: data <= 8'h00;
            16'd31446: data <= 8'h1F;
            16'd31447: data <= 8'h00;
            16'd31448: data <= 8'h1F;
            16'd31449: data <= 8'h00;
            16'd31450: data <= 8'h1F;
            16'd31451: data <= 8'h00;
            16'd31452: data <= 8'h1F;
            16'd31453: data <= 8'h00;
            16'd31454: data <= 8'h1F;
            16'd31455: data <= 8'h00;
            16'd31456: data <= 8'h1F;
            16'd31457: data <= 8'h00;
            16'd31458: data <= 8'h1F;
            16'd31459: data <= 8'h00;
            16'd31460: data <= 8'h1F;
            16'd31461: data <= 8'h00;
            16'd31462: data <= 8'h1F;
            16'd31463: data <= 8'h00;
            16'd31464: data <= 8'h1F;
            16'd31465: data <= 8'h00;
            16'd31466: data <= 8'h1F;
            16'd31467: data <= 8'h00;
            16'd31468: data <= 8'h1F;
            16'd31469: data <= 8'h00;
            16'd31470: data <= 8'h1F;
            16'd31471: data <= 8'h00;
            16'd31472: data <= 8'h1F;
            16'd31473: data <= 8'h00;
            16'd31474: data <= 8'h1F;
            16'd31475: data <= 8'h00;
            16'd31476: data <= 8'h1F;
            16'd31477: data <= 8'h00;
            16'd31478: data <= 8'h1F;
            16'd31479: data <= 8'h00;
            16'd31480: data <= 8'hFF;
            16'd31481: data <= 8'hFF;
            16'd31482: data <= 8'h1F;
            16'd31483: data <= 8'h00;
            16'd31484: data <= 8'h1F;
            16'd31485: data <= 8'h00;
            16'd31486: data <= 8'h1F;
            16'd31487: data <= 8'h00;
            16'd31488: data <= 8'h1F;
            16'd31489: data <= 8'h00;
            16'd31490: data <= 8'h1F;
            16'd31491: data <= 8'h00;
            16'd31492: data <= 8'h1F;
            16'd31493: data <= 8'h00;
            16'd31494: data <= 8'h1F;
            16'd31495: data <= 8'h00;
            16'd31496: data <= 8'h1F;
            16'd31497: data <= 8'h00;
            16'd31498: data <= 8'h1F;
            16'd31499: data <= 8'h00;
            16'd31500: data <= 8'h1F;
            16'd31501: data <= 8'h00;
            16'd31502: data <= 8'h1F;
            16'd31503: data <= 8'h00;
            16'd31504: data <= 8'h1F;
            16'd31505: data <= 8'h00;
            16'd31506: data <= 8'h1F;
            16'd31507: data <= 8'h00;
            16'd31508: data <= 8'h1F;
            16'd31509: data <= 8'h00;
            16'd31510: data <= 8'h1F;
            16'd31511: data <= 8'h00;
            16'd31512: data <= 8'h1F;
            16'd31513: data <= 8'h00;
            16'd31514: data <= 8'h1F;
            16'd31515: data <= 8'h00;
            16'd31516: data <= 8'h1F;
            16'd31517: data <= 8'h00;
            16'd31518: data <= 8'h1F;
            16'd31519: data <= 8'h00;
            16'd31520: data <= 8'hFF;
            16'd31521: data <= 8'hFF;
            16'd31522: data <= 8'h1F;
            16'd31523: data <= 8'h00;
            16'd31524: data <= 8'h1F;
            16'd31525: data <= 8'h00;
            16'd31526: data <= 8'h1F;
            16'd31527: data <= 8'h00;
            16'd31528: data <= 8'h1F;
            16'd31529: data <= 8'h00;
            16'd31530: data <= 8'h1F;
            16'd31531: data <= 8'h00;
            16'd31532: data <= 8'h1F;
            16'd31533: data <= 8'h00;
            16'd31534: data <= 8'h1F;
            16'd31535: data <= 8'h00;
            16'd31536: data <= 8'h1F;
            16'd31537: data <= 8'h00;
            16'd31538: data <= 8'h1F;
            16'd31539: data <= 8'h00;
            16'd31540: data <= 8'h1F;
            16'd31541: data <= 8'h00;
            16'd31542: data <= 8'h1F;
            16'd31543: data <= 8'h00;
            16'd31544: data <= 8'h1F;
            16'd31545: data <= 8'h00;
            16'd31546: data <= 8'h1F;
            16'd31547: data <= 8'h00;
            16'd31548: data <= 8'h1F;
            16'd31549: data <= 8'h00;
            16'd31550: data <= 8'h1F;
            16'd31551: data <= 8'h00;
            16'd31552: data <= 8'h1F;
            16'd31553: data <= 8'h00;
            16'd31554: data <= 8'h1F;
            16'd31555: data <= 8'h00;
            16'd31556: data <= 8'h1F;
            16'd31557: data <= 8'h00;
            16'd31558: data <= 8'h1F;
            16'd31559: data <= 8'h00;
            16'd31560: data <= 8'hFF;
            16'd31561: data <= 8'hFF;
            16'd31562: data <= 8'h1F;
            16'd31563: data <= 8'h00;
            16'd31564: data <= 8'h1F;
            16'd31565: data <= 8'h00;
            16'd31566: data <= 8'h1F;
            16'd31567: data <= 8'h00;
            16'd31568: data <= 8'h1F;
            16'd31569: data <= 8'h00;
            16'd31570: data <= 8'h1F;
            16'd31571: data <= 8'h00;
            16'd31572: data <= 8'h1F;
            16'd31573: data <= 8'h00;
            16'd31574: data <= 8'h1F;
            16'd31575: data <= 8'h00;
            16'd31576: data <= 8'h1F;
            16'd31577: data <= 8'h00;
            16'd31578: data <= 8'h1F;
            16'd31579: data <= 8'h00;
            16'd31580: data <= 8'h1F;
            16'd31581: data <= 8'h00;
            16'd31582: data <= 8'h1F;
            16'd31583: data <= 8'h00;
            16'd31584: data <= 8'h1F;
            16'd31585: data <= 8'h00;
            16'd31586: data <= 8'h1F;
            16'd31587: data <= 8'h00;
            16'd31588: data <= 8'h1F;
            16'd31589: data <= 8'h00;
            16'd31590: data <= 8'h1F;
            16'd31591: data <= 8'h00;
            16'd31592: data <= 8'h1F;
            16'd31593: data <= 8'h00;
            16'd31594: data <= 8'h1F;
            16'd31595: data <= 8'h00;
            16'd31596: data <= 8'h1F;
            16'd31597: data <= 8'h00;
            16'd31598: data <= 8'h1F;
            16'd31599: data <= 8'h00;
            16'd31600: data <= 8'hFF;
            16'd31601: data <= 8'hFF;
            16'd31602: data <= 8'h1F;
            16'd31603: data <= 8'h00;
            16'd31604: data <= 8'h1F;
            16'd31605: data <= 8'h00;
            16'd31606: data <= 8'h1F;
            16'd31607: data <= 8'h00;
            16'd31608: data <= 8'h1F;
            16'd31609: data <= 8'h00;
            16'd31610: data <= 8'h1F;
            16'd31611: data <= 8'h00;
            16'd31612: data <= 8'h1F;
            16'd31613: data <= 8'h00;
            16'd31614: data <= 8'h1F;
            16'd31615: data <= 8'h00;
            16'd31616: data <= 8'h1F;
            16'd31617: data <= 8'h00;
            16'd31618: data <= 8'h1F;
            16'd31619: data <= 8'h00;
            16'd31620: data <= 8'h1F;
            16'd31621: data <= 8'h00;
            16'd31622: data <= 8'h1F;
            16'd31623: data <= 8'h00;
            16'd31624: data <= 8'h1F;
            16'd31625: data <= 8'h00;
            16'd31626: data <= 8'h1F;
            16'd31627: data <= 8'h00;
            16'd31628: data <= 8'h1F;
            16'd31629: data <= 8'h00;
            16'd31630: data <= 8'h1F;
            16'd31631: data <= 8'h00;
            16'd31632: data <= 8'h1F;
            16'd31633: data <= 8'h00;
            16'd31634: data <= 8'h1F;
            16'd31635: data <= 8'h00;
            16'd31636: data <= 8'h1F;
            16'd31637: data <= 8'h00;
            16'd31638: data <= 8'h1F;
            16'd31639: data <= 8'h00;
            16'd31640: data <= 8'hFF;
            16'd31641: data <= 8'hFF;
            16'd31642: data <= 8'h1F;
            16'd31643: data <= 8'h00;
            16'd31644: data <= 8'h1F;
            16'd31645: data <= 8'h00;
            16'd31646: data <= 8'h1F;
            16'd31647: data <= 8'h00;
            16'd31648: data <= 8'h1F;
            16'd31649: data <= 8'h00;
            16'd31650: data <= 8'h1F;
            16'd31651: data <= 8'h00;
            16'd31652: data <= 8'h1F;
            16'd31653: data <= 8'h00;
            16'd31654: data <= 8'h1F;
            16'd31655: data <= 8'h00;
            16'd31656: data <= 8'h1F;
            16'd31657: data <= 8'h00;
            16'd31658: data <= 8'h1F;
            16'd31659: data <= 8'h00;
            16'd31660: data <= 8'h1F;
            16'd31661: data <= 8'h00;
            16'd31662: data <= 8'h1F;
            16'd31663: data <= 8'h00;
            16'd31664: data <= 8'h1F;
            16'd31665: data <= 8'h00;
            16'd31666: data <= 8'h1F;
            16'd31667: data <= 8'h00;
            16'd31668: data <= 8'h1F;
            16'd31669: data <= 8'h00;
            16'd31670: data <= 8'h1F;
            16'd31671: data <= 8'h00;
            16'd31672: data <= 8'h1F;
            16'd31673: data <= 8'h00;
            16'd31674: data <= 8'h1F;
            16'd31675: data <= 8'h00;
            16'd31676: data <= 8'h1F;
            16'd31677: data <= 8'h00;
            16'd31678: data <= 8'h1F;
            16'd31679: data <= 8'h00;
            16'd31680: data <= 8'hFF;
            16'd31681: data <= 8'hFF;
            16'd31682: data <= 8'h1F;
            16'd31683: data <= 8'h00;
            16'd31684: data <= 8'h1F;
            16'd31685: data <= 8'h00;
            16'd31686: data <= 8'h1F;
            16'd31687: data <= 8'h00;
            16'd31688: data <= 8'h1F;
            16'd31689: data <= 8'h00;
            16'd31690: data <= 8'h1F;
            16'd31691: data <= 8'h00;
            16'd31692: data <= 8'h1F;
            16'd31693: data <= 8'h00;
            16'd31694: data <= 8'h1F;
            16'd31695: data <= 8'h00;
            16'd31696: data <= 8'h1F;
            16'd31697: data <= 8'h00;
            16'd31698: data <= 8'h1F;
            16'd31699: data <= 8'h00;
            16'd31700: data <= 8'h1F;
            16'd31701: data <= 8'h00;
            16'd31702: data <= 8'h1F;
            16'd31703: data <= 8'h00;
            16'd31704: data <= 8'h1F;
            16'd31705: data <= 8'h00;
            16'd31706: data <= 8'h1F;
            16'd31707: data <= 8'h00;
            16'd31708: data <= 8'h1F;
            16'd31709: data <= 8'h00;
            16'd31710: data <= 8'h1F;
            16'd31711: data <= 8'h00;
            16'd31712: data <= 8'h1F;
            16'd31713: data <= 8'h00;
            16'd31714: data <= 8'h1F;
            16'd31715: data <= 8'h00;
            16'd31716: data <= 8'h1F;
            16'd31717: data <= 8'h00;
            16'd31718: data <= 8'h1F;
            16'd31719: data <= 8'h00;
            16'd31720: data <= 8'hFF;
            16'd31721: data <= 8'hFF;
            16'd31722: data <= 8'h1F;
            16'd31723: data <= 8'h00;
            16'd31724: data <= 8'h1F;
            16'd31725: data <= 8'h00;
            16'd31726: data <= 8'h1F;
            16'd31727: data <= 8'h00;
            16'd31728: data <= 8'h1F;
            16'd31729: data <= 8'h00;
            16'd31730: data <= 8'h1F;
            16'd31731: data <= 8'h00;
            16'd31732: data <= 8'h1F;
            16'd31733: data <= 8'h00;
            16'd31734: data <= 8'h1F;
            16'd31735: data <= 8'h00;
            16'd31736: data <= 8'h1F;
            16'd31737: data <= 8'h00;
            16'd31738: data <= 8'h1F;
            16'd31739: data <= 8'h00;
            16'd31740: data <= 8'h1F;
            16'd31741: data <= 8'h00;
            16'd31742: data <= 8'h1F;
            16'd31743: data <= 8'h00;
            16'd31744: data <= 8'h1F;
            16'd31745: data <= 8'h00;
            16'd31746: data <= 8'h1F;
            16'd31747: data <= 8'h00;
            16'd31748: data <= 8'h1F;
            16'd31749: data <= 8'h00;
            16'd31750: data <= 8'h1F;
            16'd31751: data <= 8'h00;
            16'd31752: data <= 8'h1F;
            16'd31753: data <= 8'h00;
            16'd31754: data <= 8'h1F;
            16'd31755: data <= 8'h00;
            16'd31756: data <= 8'h1F;
            16'd31757: data <= 8'h00;
            16'd31758: data <= 8'h1F;
            16'd31759: data <= 8'h00;
            16'd31760: data <= 8'hFF;
            16'd31761: data <= 8'hFF;
            16'd31762: data <= 8'h1F;
            16'd31763: data <= 8'h00;
            16'd31764: data <= 8'h1F;
            16'd31765: data <= 8'h00;
            16'd31766: data <= 8'h1F;
            16'd31767: data <= 8'h00;
            16'd31768: data <= 8'h1F;
            16'd31769: data <= 8'h00;
            16'd31770: data <= 8'h1F;
            16'd31771: data <= 8'h00;
            16'd31772: data <= 8'h1F;
            16'd31773: data <= 8'h00;
            16'd31774: data <= 8'h1F;
            16'd31775: data <= 8'h00;
            16'd31776: data <= 8'h1F;
            16'd31777: data <= 8'h00;
            16'd31778: data <= 8'h1F;
            16'd31779: data <= 8'h00;
            16'd31780: data <= 8'h1F;
            16'd31781: data <= 8'h00;
            16'd31782: data <= 8'h1F;
            16'd31783: data <= 8'h00;
            16'd31784: data <= 8'h1F;
            16'd31785: data <= 8'h00;
            16'd31786: data <= 8'h1F;
            16'd31787: data <= 8'h00;
            16'd31788: data <= 8'h1F;
            16'd31789: data <= 8'h00;
            16'd31790: data <= 8'h1F;
            16'd31791: data <= 8'h00;
            16'd31792: data <= 8'h1F;
            16'd31793: data <= 8'h00;
            16'd31794: data <= 8'h1F;
            16'd31795: data <= 8'h00;
            16'd31796: data <= 8'h1F;
            16'd31797: data <= 8'h00;
            16'd31798: data <= 8'h1F;
            16'd31799: data <= 8'h00;
            16'd31800: data <= 8'hFF;
            16'd31801: data <= 8'hFF;
            16'd31802: data <= 8'h1F;
            16'd31803: data <= 8'h00;
            16'd31804: data <= 8'h1F;
            16'd31805: data <= 8'h00;
            16'd31806: data <= 8'h1F;
            16'd31807: data <= 8'h00;
            16'd31808: data <= 8'h1F;
            16'd31809: data <= 8'h00;
            16'd31810: data <= 8'h1F;
            16'd31811: data <= 8'h00;
            16'd31812: data <= 8'h1F;
            16'd31813: data <= 8'h00;
            16'd31814: data <= 8'h1F;
            16'd31815: data <= 8'h00;
            16'd31816: data <= 8'h1F;
            16'd31817: data <= 8'h00;
            16'd31818: data <= 8'h1F;
            16'd31819: data <= 8'h00;
            16'd31820: data <= 8'h1F;
            16'd31821: data <= 8'h00;
            16'd31822: data <= 8'h1F;
            16'd31823: data <= 8'h00;
            16'd31824: data <= 8'h1F;
            16'd31825: data <= 8'h00;
            16'd31826: data <= 8'h1F;
            16'd31827: data <= 8'h00;
            16'd31828: data <= 8'h1F;
            16'd31829: data <= 8'h00;
            16'd31830: data <= 8'h1F;
            16'd31831: data <= 8'h00;
            16'd31832: data <= 8'h1F;
            16'd31833: data <= 8'h00;
            16'd31834: data <= 8'h1F;
            16'd31835: data <= 8'h00;
            16'd31836: data <= 8'h1F;
            16'd31837: data <= 8'h00;
            16'd31838: data <= 8'h1F;
            16'd31839: data <= 8'h00;
            16'd31840: data <= 8'hFF;
            16'd31841: data <= 8'hFF;
            16'd31842: data <= 8'h1F;
            16'd31843: data <= 8'h00;
            16'd31844: data <= 8'h1F;
            16'd31845: data <= 8'h00;
            16'd31846: data <= 8'h1F;
            16'd31847: data <= 8'h00;
            16'd31848: data <= 8'h1F;
            16'd31849: data <= 8'h00;
            16'd31850: data <= 8'h1F;
            16'd31851: data <= 8'h00;
            16'd31852: data <= 8'h1F;
            16'd31853: data <= 8'h00;
            16'd31854: data <= 8'h1F;
            16'd31855: data <= 8'h00;
            16'd31856: data <= 8'h1F;
            16'd31857: data <= 8'h00;
            16'd31858: data <= 8'h1F;
            16'd31859: data <= 8'h00;
            16'd31860: data <= 8'h1F;
            16'd31861: data <= 8'h00;
            16'd31862: data <= 8'h1F;
            16'd31863: data <= 8'h00;
            16'd31864: data <= 8'h1F;
            16'd31865: data <= 8'h00;
            16'd31866: data <= 8'h1F;
            16'd31867: data <= 8'h00;
            16'd31868: data <= 8'h1F;
            16'd31869: data <= 8'h00;
            16'd31870: data <= 8'h1F;
            16'd31871: data <= 8'h00;
            16'd31872: data <= 8'h1F;
            16'd31873: data <= 8'h00;
            16'd31874: data <= 8'h1F;
            16'd31875: data <= 8'h00;
            16'd31876: data <= 8'h1F;
            16'd31877: data <= 8'h00;
            16'd31878: data <= 8'h1F;
            16'd31879: data <= 8'h00;
            16'd31880: data <= 8'hFF;
            16'd31881: data <= 8'hFF;
            16'd31882: data <= 8'h1F;
            16'd31883: data <= 8'h00;
            16'd31884: data <= 8'h1F;
            16'd31885: data <= 8'h00;
            16'd31886: data <= 8'h1F;
            16'd31887: data <= 8'h00;
            16'd31888: data <= 8'h1F;
            16'd31889: data <= 8'h00;
            16'd31890: data <= 8'h1F;
            16'd31891: data <= 8'h00;
            16'd31892: data <= 8'h1F;
            16'd31893: data <= 8'h00;
            16'd31894: data <= 8'h1F;
            16'd31895: data <= 8'h00;
            16'd31896: data <= 8'h1F;
            16'd31897: data <= 8'h00;
            16'd31898: data <= 8'h1F;
            16'd31899: data <= 8'h00;
            16'd31900: data <= 8'h1F;
            16'd31901: data <= 8'h00;
            16'd31902: data <= 8'h1F;
            16'd31903: data <= 8'h00;
            16'd31904: data <= 8'h1F;
            16'd31905: data <= 8'h00;
            16'd31906: data <= 8'h1F;
            16'd31907: data <= 8'h00;
            16'd31908: data <= 8'h1F;
            16'd31909: data <= 8'h00;
            16'd31910: data <= 8'h1F;
            16'd31911: data <= 8'h00;
            16'd31912: data <= 8'h1F;
            16'd31913: data <= 8'h00;
            16'd31914: data <= 8'h1F;
            16'd31915: data <= 8'h00;
            16'd31916: data <= 8'h1F;
            16'd31917: data <= 8'h00;
            16'd31918: data <= 8'h1F;
            16'd31919: data <= 8'h00;
            16'd31920: data <= 8'hFF;
            16'd31921: data <= 8'hFF;
            16'd31922: data <= 8'h1F;
            16'd31923: data <= 8'h00;
            16'd31924: data <= 8'h1F;
            16'd31925: data <= 8'h00;
            16'd31926: data <= 8'h1F;
            16'd31927: data <= 8'h00;
            16'd31928: data <= 8'h1F;
            16'd31929: data <= 8'h00;
            16'd31930: data <= 8'h1F;
            16'd31931: data <= 8'h00;
            16'd31932: data <= 8'h1F;
            16'd31933: data <= 8'h00;
            16'd31934: data <= 8'h1F;
            16'd31935: data <= 8'h00;
            16'd31936: data <= 8'h1F;
            16'd31937: data <= 8'h00;
            16'd31938: data <= 8'h1F;
            16'd31939: data <= 8'h00;
            16'd31940: data <= 8'h1F;
            16'd31941: data <= 8'h00;
            16'd31942: data <= 8'h1F;
            16'd31943: data <= 8'h00;
            16'd31944: data <= 8'h1F;
            16'd31945: data <= 8'h00;
            16'd31946: data <= 8'h1F;
            16'd31947: data <= 8'h00;
            16'd31948: data <= 8'h1F;
            16'd31949: data <= 8'h00;
            16'd31950: data <= 8'h1F;
            16'd31951: data <= 8'h00;
            16'd31952: data <= 8'h1F;
            16'd31953: data <= 8'h00;
            16'd31954: data <= 8'h1F;
            16'd31955: data <= 8'h00;
            16'd31956: data <= 8'h1F;
            16'd31957: data <= 8'h00;
            16'd31958: data <= 8'h1F;
            16'd31959: data <= 8'h00;
            16'd31960: data <= 8'hFF;
            16'd31961: data <= 8'hFF;
            16'd31962: data <= 8'h1F;
            16'd31963: data <= 8'h00;
            16'd31964: data <= 8'h1F;
            16'd31965: data <= 8'h00;
            16'd31966: data <= 8'h1F;
            16'd31967: data <= 8'h00;
            16'd31968: data <= 8'h1F;
            16'd31969: data <= 8'h00;
            16'd31970: data <= 8'h1F;
            16'd31971: data <= 8'h00;
            16'd31972: data <= 8'h1F;
            16'd31973: data <= 8'h00;
            16'd31974: data <= 8'h1F;
            16'd31975: data <= 8'h00;
            16'd31976: data <= 8'h1F;
            16'd31977: data <= 8'h00;
            16'd31978: data <= 8'h1F;
            16'd31979: data <= 8'h00;
            16'd31980: data <= 8'h1F;
            16'd31981: data <= 8'h00;
            16'd31982: data <= 8'h1F;
            16'd31983: data <= 8'h00;
            16'd31984: data <= 8'h1F;
            16'd31985: data <= 8'h00;
            16'd31986: data <= 8'h1F;
            16'd31987: data <= 8'h00;
            16'd31988: data <= 8'h1F;
            16'd31989: data <= 8'h00;
            16'd31990: data <= 8'h1F;
            16'd31991: data <= 8'h00;
            16'd31992: data <= 8'h1F;
            16'd31993: data <= 8'h00;
            16'd31994: data <= 8'h1F;
            16'd31995: data <= 8'h00;
            16'd31996: data <= 8'h1F;
            16'd31997: data <= 8'h00;
            16'd31998: data <= 8'h1F;
            16'd31999: data <= 8'h00;
            16'd32000: data <= 8'hFF;
            16'd32001: data <= 8'hFF;
            16'd32002: data <= 8'h1F;
            16'd32003: data <= 8'h00;
            16'd32004: data <= 8'h1F;
            16'd32005: data <= 8'h00;
            16'd32006: data <= 8'h1F;
            16'd32007: data <= 8'h00;
            16'd32008: data <= 8'h1F;
            16'd32009: data <= 8'h00;
            16'd32010: data <= 8'h1F;
            16'd32011: data <= 8'h00;
            16'd32012: data <= 8'h1F;
            16'd32013: data <= 8'h00;
            16'd32014: data <= 8'h1F;
            16'd32015: data <= 8'h00;
            16'd32016: data <= 8'h1F;
            16'd32017: data <= 8'h00;
            16'd32018: data <= 8'h1F;
            16'd32019: data <= 8'h00;
            16'd32020: data <= 8'h1F;
            16'd32021: data <= 8'h00;
            16'd32022: data <= 8'h1F;
            16'd32023: data <= 8'h00;
            16'd32024: data <= 8'h1F;
            16'd32025: data <= 8'h00;
            16'd32026: data <= 8'h1F;
            16'd32027: data <= 8'h00;
            16'd32028: data <= 8'h1F;
            16'd32029: data <= 8'h00;
            16'd32030: data <= 8'h1F;
            16'd32031: data <= 8'h00;
            16'd32032: data <= 8'h1F;
            16'd32033: data <= 8'h00;
            16'd32034: data <= 8'h1F;
            16'd32035: data <= 8'h00;
            16'd32036: data <= 8'h1F;
            16'd32037: data <= 8'h00;
            16'd32038: data <= 8'h1F;
            16'd32039: data <= 8'h00;
            16'd32040: data <= 8'hFF;
            16'd32041: data <= 8'hFF;
            16'd32042: data <= 8'h1F;
            16'd32043: data <= 8'h00;
            16'd32044: data <= 8'h1F;
            16'd32045: data <= 8'h00;
            16'd32046: data <= 8'h1F;
            16'd32047: data <= 8'h00;
            16'd32048: data <= 8'h1F;
            16'd32049: data <= 8'h00;
            16'd32050: data <= 8'h1F;
            16'd32051: data <= 8'h00;
            16'd32052: data <= 8'h1F;
            16'd32053: data <= 8'h00;
            16'd32054: data <= 8'h1F;
            16'd32055: data <= 8'h00;
            16'd32056: data <= 8'h1F;
            16'd32057: data <= 8'h00;
            16'd32058: data <= 8'h1F;
            16'd32059: data <= 8'h00;
            16'd32060: data <= 8'h1F;
            16'd32061: data <= 8'h00;
            16'd32062: data <= 8'h1F;
            16'd32063: data <= 8'h00;
            16'd32064: data <= 8'h1F;
            16'd32065: data <= 8'h00;
            16'd32066: data <= 8'h1F;
            16'd32067: data <= 8'h00;
            16'd32068: data <= 8'h1F;
            16'd32069: data <= 8'h00;
            16'd32070: data <= 8'h1F;
            16'd32071: data <= 8'h00;
            16'd32072: data <= 8'h1F;
            16'd32073: data <= 8'h00;
            16'd32074: data <= 8'h1F;
            16'd32075: data <= 8'h00;
            16'd32076: data <= 8'h1F;
            16'd32077: data <= 8'h00;
            16'd32078: data <= 8'h1F;
            16'd32079: data <= 8'h00;
            16'd32080: data <= 8'hFF;
            16'd32081: data <= 8'hFF;
            16'd32082: data <= 8'h1F;
            16'd32083: data <= 8'h00;
            16'd32084: data <= 8'h1F;
            16'd32085: data <= 8'h00;
            16'd32086: data <= 8'h1F;
            16'd32087: data <= 8'h00;
            16'd32088: data <= 8'h1F;
            16'd32089: data <= 8'h00;
            16'd32090: data <= 8'h1F;
            16'd32091: data <= 8'h00;
            16'd32092: data <= 8'h1F;
            16'd32093: data <= 8'h00;
            16'd32094: data <= 8'h1F;
            16'd32095: data <= 8'h00;
            16'd32096: data <= 8'h1F;
            16'd32097: data <= 8'h00;
            16'd32098: data <= 8'h1F;
            16'd32099: data <= 8'h00;
            16'd32100: data <= 8'h1F;
            16'd32101: data <= 8'h00;
            16'd32102: data <= 8'h1F;
            16'd32103: data <= 8'h00;
            16'd32104: data <= 8'h1F;
            16'd32105: data <= 8'h00;
            16'd32106: data <= 8'h1F;
            16'd32107: data <= 8'h00;
            16'd32108: data <= 8'h1F;
            16'd32109: data <= 8'h00;
            16'd32110: data <= 8'h1F;
            16'd32111: data <= 8'h00;
            16'd32112: data <= 8'h1F;
            16'd32113: data <= 8'h00;
            16'd32114: data <= 8'h1F;
            16'd32115: data <= 8'h00;
            16'd32116: data <= 8'h1F;
            16'd32117: data <= 8'h00;
            16'd32118: data <= 8'h1F;
            16'd32119: data <= 8'h00;
            16'd32120: data <= 8'hFF;
            16'd32121: data <= 8'hFF;
            16'd32122: data <= 8'h1F;
            16'd32123: data <= 8'h00;
            16'd32124: data <= 8'h1F;
            16'd32125: data <= 8'h00;
            16'd32126: data <= 8'h1F;
            16'd32127: data <= 8'h00;
            16'd32128: data <= 8'h1F;
            16'd32129: data <= 8'h00;
            16'd32130: data <= 8'h1F;
            16'd32131: data <= 8'h00;
            16'd32132: data <= 8'h1F;
            16'd32133: data <= 8'h00;
            16'd32134: data <= 8'h1F;
            16'd32135: data <= 8'h00;
            16'd32136: data <= 8'h1F;
            16'd32137: data <= 8'h00;
            16'd32138: data <= 8'h1F;
            16'd32139: data <= 8'h00;
            16'd32140: data <= 8'h1F;
            16'd32141: data <= 8'h00;
            16'd32142: data <= 8'h1F;
            16'd32143: data <= 8'h00;
            16'd32144: data <= 8'h1F;
            16'd32145: data <= 8'h00;
            16'd32146: data <= 8'h1F;
            16'd32147: data <= 8'h00;
            16'd32148: data <= 8'h1F;
            16'd32149: data <= 8'h00;
            16'd32150: data <= 8'h1F;
            16'd32151: data <= 8'h00;
            16'd32152: data <= 8'h1F;
            16'd32153: data <= 8'h00;
            16'd32154: data <= 8'h1F;
            16'd32155: data <= 8'h00;
            16'd32156: data <= 8'h1F;
            16'd32157: data <= 8'h00;
            16'd32158: data <= 8'h1F;
            16'd32159: data <= 8'h00;
            16'd32160: data <= 8'hFF;
            16'd32161: data <= 8'hFF;
            16'd32162: data <= 8'h1F;
            16'd32163: data <= 8'h00;
            16'd32164: data <= 8'h1F;
            16'd32165: data <= 8'h00;
            16'd32166: data <= 8'h1F;
            16'd32167: data <= 8'h00;
            16'd32168: data <= 8'h1F;
            16'd32169: data <= 8'h00;
            16'd32170: data <= 8'h1F;
            16'd32171: data <= 8'h00;
            16'd32172: data <= 8'h1F;
            16'd32173: data <= 8'h00;
            16'd32174: data <= 8'h1F;
            16'd32175: data <= 8'h00;
            16'd32176: data <= 8'h1F;
            16'd32177: data <= 8'h00;
            16'd32178: data <= 8'h1F;
            16'd32179: data <= 8'h00;
            16'd32180: data <= 8'h1F;
            16'd32181: data <= 8'h00;
            16'd32182: data <= 8'h1F;
            16'd32183: data <= 8'h00;
            16'd32184: data <= 8'h1F;
            16'd32185: data <= 8'h00;
            16'd32186: data <= 8'h1F;
            16'd32187: data <= 8'h00;
            16'd32188: data <= 8'h1F;
            16'd32189: data <= 8'h00;
            16'd32190: data <= 8'h1F;
            16'd32191: data <= 8'h00;
            16'd32192: data <= 8'h1F;
            16'd32193: data <= 8'h00;
            16'd32194: data <= 8'h1F;
            16'd32195: data <= 8'h00;
            16'd32196: data <= 8'h1F;
            16'd32197: data <= 8'h00;
            16'd32198: data <= 8'h1F;
            16'd32199: data <= 8'h00;
            16'd32200: data <= 8'hFF;
            16'd32201: data <= 8'hFF;
            16'd32202: data <= 8'h1F;
            16'd32203: data <= 8'h00;
            16'd32204: data <= 8'h1F;
            16'd32205: data <= 8'h00;
            16'd32206: data <= 8'h1F;
            16'd32207: data <= 8'h00;
            16'd32208: data <= 8'h1F;
            16'd32209: data <= 8'h00;
            16'd32210: data <= 8'h1F;
            16'd32211: data <= 8'h00;
            16'd32212: data <= 8'h1F;
            16'd32213: data <= 8'h00;
            16'd32214: data <= 8'h1F;
            16'd32215: data <= 8'h00;
            16'd32216: data <= 8'h1F;
            16'd32217: data <= 8'h00;
            16'd32218: data <= 8'h1F;
            16'd32219: data <= 8'h00;
            16'd32220: data <= 8'h1F;
            16'd32221: data <= 8'h00;
            16'd32222: data <= 8'h1F;
            16'd32223: data <= 8'h00;
            16'd32224: data <= 8'h1F;
            16'd32225: data <= 8'h00;
            16'd32226: data <= 8'h1F;
            16'd32227: data <= 8'h00;
            16'd32228: data <= 8'h1F;
            16'd32229: data <= 8'h00;
            16'd32230: data <= 8'h1F;
            16'd32231: data <= 8'h00;
            16'd32232: data <= 8'h1F;
            16'd32233: data <= 8'h00;
            16'd32234: data <= 8'h1F;
            16'd32235: data <= 8'h00;
            16'd32236: data <= 8'h1F;
            16'd32237: data <= 8'h00;
            16'd32238: data <= 8'h1F;
            16'd32239: data <= 8'h00;
            16'd32240: data <= 8'hFF;
            16'd32241: data <= 8'hFF;
            16'd32242: data <= 8'h1F;
            16'd32243: data <= 8'h00;
            16'd32244: data <= 8'h1F;
            16'd32245: data <= 8'h00;
            16'd32246: data <= 8'h1F;
            16'd32247: data <= 8'h00;
            16'd32248: data <= 8'h1F;
            16'd32249: data <= 8'h00;
            16'd32250: data <= 8'h1F;
            16'd32251: data <= 8'h00;
            16'd32252: data <= 8'h1F;
            16'd32253: data <= 8'h00;
            16'd32254: data <= 8'h1F;
            16'd32255: data <= 8'h00;
            16'd32256: data <= 8'h1F;
            16'd32257: data <= 8'h00;
            16'd32258: data <= 8'h1F;
            16'd32259: data <= 8'h00;
            16'd32260: data <= 8'h1F;
            16'd32261: data <= 8'h00;
            16'd32262: data <= 8'h1F;
            16'd32263: data <= 8'h00;
            16'd32264: data <= 8'h1F;
            16'd32265: data <= 8'h00;
            16'd32266: data <= 8'h1F;
            16'd32267: data <= 8'h00;
            16'd32268: data <= 8'h1F;
            16'd32269: data <= 8'h00;
            16'd32270: data <= 8'h1F;
            16'd32271: data <= 8'h00;
            16'd32272: data <= 8'h1F;
            16'd32273: data <= 8'h00;
            16'd32274: data <= 8'h1F;
            16'd32275: data <= 8'h00;
            16'd32276: data <= 8'h1F;
            16'd32277: data <= 8'h00;
            16'd32278: data <= 8'h1F;
            16'd32279: data <= 8'h00;
            16'd32280: data <= 8'hFF;
            16'd32281: data <= 8'hFF;
            16'd32282: data <= 8'h1F;
            16'd32283: data <= 8'h00;
            16'd32284: data <= 8'h1F;
            16'd32285: data <= 8'h00;
            16'd32286: data <= 8'h1F;
            16'd32287: data <= 8'h00;
            16'd32288: data <= 8'h1F;
            16'd32289: data <= 8'h00;
            16'd32290: data <= 8'h1F;
            16'd32291: data <= 8'h00;
            16'd32292: data <= 8'h1F;
            16'd32293: data <= 8'h00;
            16'd32294: data <= 8'h1F;
            16'd32295: data <= 8'h00;
            16'd32296: data <= 8'h1F;
            16'd32297: data <= 8'h00;
            16'd32298: data <= 8'h1F;
            16'd32299: data <= 8'h00;
            16'd32300: data <= 8'h1F;
            16'd32301: data <= 8'h00;
            16'd32302: data <= 8'h1F;
            16'd32303: data <= 8'h00;
            16'd32304: data <= 8'h1F;
            16'd32305: data <= 8'h00;
            16'd32306: data <= 8'h1F;
            16'd32307: data <= 8'h00;
            16'd32308: data <= 8'h1F;
            16'd32309: data <= 8'h00;
            16'd32310: data <= 8'h1F;
            16'd32311: data <= 8'h00;
            16'd32312: data <= 8'h1F;
            16'd32313: data <= 8'h00;
            16'd32314: data <= 8'h1F;
            16'd32315: data <= 8'h00;
            16'd32316: data <= 8'h1F;
            16'd32317: data <= 8'h00;
            16'd32318: data <= 8'h1F;
            16'd32319: data <= 8'h00;
            16'd32320: data <= 8'hFF;
            16'd32321: data <= 8'hFF;
            16'd32322: data <= 8'h1F;
            16'd32323: data <= 8'h00;
            16'd32324: data <= 8'h1F;
            16'd32325: data <= 8'h00;
            16'd32326: data <= 8'h1F;
            16'd32327: data <= 8'h00;
            16'd32328: data <= 8'h1F;
            16'd32329: data <= 8'h00;
            16'd32330: data <= 8'h1F;
            16'd32331: data <= 8'h00;
            16'd32332: data <= 8'h1F;
            16'd32333: data <= 8'h00;
            16'd32334: data <= 8'h1F;
            16'd32335: data <= 8'h00;
            16'd32336: data <= 8'h1F;
            16'd32337: data <= 8'h00;
            16'd32338: data <= 8'h1F;
            16'd32339: data <= 8'h00;
            16'd32340: data <= 8'h1F;
            16'd32341: data <= 8'h00;
            16'd32342: data <= 8'h1F;
            16'd32343: data <= 8'h00;
            16'd32344: data <= 8'h1F;
            16'd32345: data <= 8'h00;
            16'd32346: data <= 8'h1F;
            16'd32347: data <= 8'h00;
            16'd32348: data <= 8'h1F;
            16'd32349: data <= 8'h00;
            16'd32350: data <= 8'h1F;
            16'd32351: data <= 8'h00;
            16'd32352: data <= 8'h1F;
            16'd32353: data <= 8'h00;
            16'd32354: data <= 8'h1F;
            16'd32355: data <= 8'h00;
            16'd32356: data <= 8'h1F;
            16'd32357: data <= 8'h00;
            16'd32358: data <= 8'h1F;
            16'd32359: data <= 8'h00;
            16'd32360: data <= 8'hFF;
            16'd32361: data <= 8'hFF;
            16'd32362: data <= 8'h1F;
            16'd32363: data <= 8'h00;
            16'd32364: data <= 8'h1F;
            16'd32365: data <= 8'h00;
            16'd32366: data <= 8'h1F;
            16'd32367: data <= 8'h00;
            16'd32368: data <= 8'h1F;
            16'd32369: data <= 8'h00;
            16'd32370: data <= 8'h1F;
            16'd32371: data <= 8'h00;
            16'd32372: data <= 8'h1F;
            16'd32373: data <= 8'h00;
            16'd32374: data <= 8'h1F;
            16'd32375: data <= 8'h00;
            16'd32376: data <= 8'h1F;
            16'd32377: data <= 8'h00;
            16'd32378: data <= 8'h1F;
            16'd32379: data <= 8'h00;
            16'd32380: data <= 8'h1F;
            16'd32381: data <= 8'h00;
            16'd32382: data <= 8'h1F;
            16'd32383: data <= 8'h00;
            16'd32384: data <= 8'h1F;
            16'd32385: data <= 8'h00;
            16'd32386: data <= 8'h1F;
            16'd32387: data <= 8'h00;
            16'd32388: data <= 8'h1F;
            16'd32389: data <= 8'h00;
            16'd32390: data <= 8'h1F;
            16'd32391: data <= 8'h00;
            16'd32392: data <= 8'h1F;
            16'd32393: data <= 8'h00;
            16'd32394: data <= 8'h1F;
            16'd32395: data <= 8'h00;
            16'd32396: data <= 8'h1F;
            16'd32397: data <= 8'h00;
            16'd32398: data <= 8'h1F;
            16'd32399: data <= 8'h00;
            16'd32400: data <= 8'hFF;
            16'd32401: data <= 8'hFF;
            16'd32402: data <= 8'h1F;
            16'd32403: data <= 8'h00;
            16'd32404: data <= 8'h1F;
            16'd32405: data <= 8'h00;
            16'd32406: data <= 8'h1F;
            16'd32407: data <= 8'h00;
            16'd32408: data <= 8'h1F;
            16'd32409: data <= 8'h00;
            16'd32410: data <= 8'h1F;
            16'd32411: data <= 8'h00;
            16'd32412: data <= 8'h1F;
            16'd32413: data <= 8'h00;
            16'd32414: data <= 8'h1F;
            16'd32415: data <= 8'h00;
            16'd32416: data <= 8'h1F;
            16'd32417: data <= 8'h00;
            16'd32418: data <= 8'h1F;
            16'd32419: data <= 8'h00;
            16'd32420: data <= 8'h1F;
            16'd32421: data <= 8'h00;
            16'd32422: data <= 8'h1F;
            16'd32423: data <= 8'h00;
            16'd32424: data <= 8'h1F;
            16'd32425: data <= 8'h00;
            16'd32426: data <= 8'h1F;
            16'd32427: data <= 8'h00;
            16'd32428: data <= 8'h1F;
            16'd32429: data <= 8'h00;
            16'd32430: data <= 8'h1F;
            16'd32431: data <= 8'h00;
            16'd32432: data <= 8'h1F;
            16'd32433: data <= 8'h00;
            16'd32434: data <= 8'h1F;
            16'd32435: data <= 8'h00;
            16'd32436: data <= 8'h1F;
            16'd32437: data <= 8'h00;
            16'd32438: data <= 8'h1F;
            16'd32439: data <= 8'h00;
            16'd32440: data <= 8'hFF;
            16'd32441: data <= 8'hFF;
            16'd32442: data <= 8'h1F;
            16'd32443: data <= 8'h00;
            16'd32444: data <= 8'h1F;
            16'd32445: data <= 8'h00;
            16'd32446: data <= 8'h1F;
            16'd32447: data <= 8'h00;
            16'd32448: data <= 8'h1F;
            16'd32449: data <= 8'h00;
            16'd32450: data <= 8'h1F;
            16'd32451: data <= 8'h00;
            16'd32452: data <= 8'h1F;
            16'd32453: data <= 8'h00;
            16'd32454: data <= 8'h1F;
            16'd32455: data <= 8'h00;
            16'd32456: data <= 8'h1F;
            16'd32457: data <= 8'h00;
            16'd32458: data <= 8'h1F;
            16'd32459: data <= 8'h00;
            16'd32460: data <= 8'h1F;
            16'd32461: data <= 8'h00;
            16'd32462: data <= 8'h1F;
            16'd32463: data <= 8'h00;
            16'd32464: data <= 8'h1F;
            16'd32465: data <= 8'h00;
            16'd32466: data <= 8'h1F;
            16'd32467: data <= 8'h00;
            16'd32468: data <= 8'h1F;
            16'd32469: data <= 8'h00;
            16'd32470: data <= 8'h1F;
            16'd32471: data <= 8'h00;
            16'd32472: data <= 8'h1F;
            16'd32473: data <= 8'h00;
            16'd32474: data <= 8'h1F;
            16'd32475: data <= 8'h00;
            16'd32476: data <= 8'h1F;
            16'd32477: data <= 8'h00;
            16'd32478: data <= 8'h1F;
            16'd32479: data <= 8'h00;
            16'd32480: data <= 8'hFF;
            16'd32481: data <= 8'hFF;
            16'd32482: data <= 8'h1F;
            16'd32483: data <= 8'h00;
            16'd32484: data <= 8'h1F;
            16'd32485: data <= 8'h00;
            16'd32486: data <= 8'h1F;
            16'd32487: data <= 8'h00;
            16'd32488: data <= 8'h1F;
            16'd32489: data <= 8'h00;
            16'd32490: data <= 8'h1F;
            16'd32491: data <= 8'h00;
            16'd32492: data <= 8'h1F;
            16'd32493: data <= 8'h00;
            16'd32494: data <= 8'h1F;
            16'd32495: data <= 8'h00;
            16'd32496: data <= 8'h1F;
            16'd32497: data <= 8'h00;
            16'd32498: data <= 8'h1F;
            16'd32499: data <= 8'h00;
            16'd32500: data <= 8'h1F;
            16'd32501: data <= 8'h00;
            16'd32502: data <= 8'h1F;
            16'd32503: data <= 8'h00;
            16'd32504: data <= 8'h1F;
            16'd32505: data <= 8'h00;
            16'd32506: data <= 8'h1F;
            16'd32507: data <= 8'h00;
            16'd32508: data <= 8'h1F;
            16'd32509: data <= 8'h00;
            16'd32510: data <= 8'h1F;
            16'd32511: data <= 8'h00;
            16'd32512: data <= 8'h1F;
            16'd32513: data <= 8'h00;
            16'd32514: data <= 8'h1F;
            16'd32515: data <= 8'h00;
            16'd32516: data <= 8'h1F;
            16'd32517: data <= 8'h00;
            16'd32518: data <= 8'h1F;
            16'd32519: data <= 8'h00;
            16'd32520: data <= 8'hFF;
            16'd32521: data <= 8'hFF;
            16'd32522: data <= 8'h1F;
            16'd32523: data <= 8'h00;
            16'd32524: data <= 8'h1F;
            16'd32525: data <= 8'h00;
            16'd32526: data <= 8'h1F;
            16'd32527: data <= 8'h00;
            16'd32528: data <= 8'h1F;
            16'd32529: data <= 8'h00;
            16'd32530: data <= 8'h1F;
            16'd32531: data <= 8'h00;
            16'd32532: data <= 8'h1F;
            16'd32533: data <= 8'h00;
            16'd32534: data <= 8'h1F;
            16'd32535: data <= 8'h00;
            16'd32536: data <= 8'h1F;
            16'd32537: data <= 8'h00;
            16'd32538: data <= 8'h1F;
            16'd32539: data <= 8'h00;
            16'd32540: data <= 8'h1F;
            16'd32541: data <= 8'h00;
            16'd32542: data <= 8'h1F;
            16'd32543: data <= 8'h00;
            16'd32544: data <= 8'h1F;
            16'd32545: data <= 8'h00;
            16'd32546: data <= 8'h1F;
            16'd32547: data <= 8'h00;
            16'd32548: data <= 8'h1F;
            16'd32549: data <= 8'h00;
            16'd32550: data <= 8'h1F;
            16'd32551: data <= 8'h00;
            16'd32552: data <= 8'h1F;
            16'd32553: data <= 8'h00;
            16'd32554: data <= 8'h1F;
            16'd32555: data <= 8'h00;
            16'd32556: data <= 8'h1F;
            16'd32557: data <= 8'h00;
            16'd32558: data <= 8'h1F;
            16'd32559: data <= 8'h00;
            16'd32560: data <= 8'hFF;
            16'd32561: data <= 8'hFF;
            16'd32562: data <= 8'h1F;
            16'd32563: data <= 8'h00;
            16'd32564: data <= 8'h1F;
            16'd32565: data <= 8'h00;
            16'd32566: data <= 8'h1F;
            16'd32567: data <= 8'h00;
            16'd32568: data <= 8'h1F;
            16'd32569: data <= 8'h00;
            16'd32570: data <= 8'h1F;
            16'd32571: data <= 8'h00;
            16'd32572: data <= 8'h1F;
            16'd32573: data <= 8'h00;
            16'd32574: data <= 8'h1F;
            16'd32575: data <= 8'h00;
            16'd32576: data <= 8'h1F;
            16'd32577: data <= 8'h00;
            16'd32578: data <= 8'h1F;
            16'd32579: data <= 8'h00;
            16'd32580: data <= 8'h1F;
            16'd32581: data <= 8'h00;
            16'd32582: data <= 8'h1F;
            16'd32583: data <= 8'h00;
            16'd32584: data <= 8'h1F;
            16'd32585: data <= 8'h00;
            16'd32586: data <= 8'h1F;
            16'd32587: data <= 8'h00;
            16'd32588: data <= 8'h1F;
            16'd32589: data <= 8'h00;
            16'd32590: data <= 8'h1F;
            16'd32591: data <= 8'h00;
            16'd32592: data <= 8'h1F;
            16'd32593: data <= 8'h00;
            16'd32594: data <= 8'h1F;
            16'd32595: data <= 8'h00;
            16'd32596: data <= 8'h1F;
            16'd32597: data <= 8'h00;
            16'd32598: data <= 8'h1F;
            16'd32599: data <= 8'h00;
            16'd32600: data <= 8'hFF;
            16'd32601: data <= 8'hFF;
            16'd32602: data <= 8'h1F;
            16'd32603: data <= 8'h00;
            16'd32604: data <= 8'h1F;
            16'd32605: data <= 8'h00;
            16'd32606: data <= 8'h1F;
            16'd32607: data <= 8'h00;
            16'd32608: data <= 8'h1F;
            16'd32609: data <= 8'h00;
            16'd32610: data <= 8'h1F;
            16'd32611: data <= 8'h00;
            16'd32612: data <= 8'h1F;
            16'd32613: data <= 8'h00;
            16'd32614: data <= 8'h1F;
            16'd32615: data <= 8'h00;
            16'd32616: data <= 8'h1F;
            16'd32617: data <= 8'h00;
            16'd32618: data <= 8'h1F;
            16'd32619: data <= 8'h00;
            16'd32620: data <= 8'h1F;
            16'd32621: data <= 8'h00;
            16'd32622: data <= 8'h1F;
            16'd32623: data <= 8'h00;
            16'd32624: data <= 8'h1F;
            16'd32625: data <= 8'h00;
            16'd32626: data <= 8'h1F;
            16'd32627: data <= 8'h00;
            16'd32628: data <= 8'h1F;
            16'd32629: data <= 8'h00;
            16'd32630: data <= 8'h1F;
            16'd32631: data <= 8'h00;
            16'd32632: data <= 8'h1F;
            16'd32633: data <= 8'h00;
            16'd32634: data <= 8'h1F;
            16'd32635: data <= 8'h00;
            16'd32636: data <= 8'h1F;
            16'd32637: data <= 8'h00;
            16'd32638: data <= 8'h1F;
            16'd32639: data <= 8'h00;
            16'd32640: data <= 8'hFF;
            16'd32641: data <= 8'hFF;
            16'd32642: data <= 8'h1F;
            16'd32643: data <= 8'h00;
            16'd32644: data <= 8'h1F;
            16'd32645: data <= 8'h00;
            16'd32646: data <= 8'h1F;
            16'd32647: data <= 8'h00;
            16'd32648: data <= 8'h1F;
            16'd32649: data <= 8'h00;
            16'd32650: data <= 8'h1F;
            16'd32651: data <= 8'h00;
            16'd32652: data <= 8'h1F;
            16'd32653: data <= 8'h00;
            16'd32654: data <= 8'h1F;
            16'd32655: data <= 8'h00;
            16'd32656: data <= 8'h1F;
            16'd32657: data <= 8'h00;
            16'd32658: data <= 8'h1F;
            16'd32659: data <= 8'h00;
            16'd32660: data <= 8'h1F;
            16'd32661: data <= 8'h00;
            16'd32662: data <= 8'h1F;
            16'd32663: data <= 8'h00;
            16'd32664: data <= 8'h1F;
            16'd32665: data <= 8'h00;
            16'd32666: data <= 8'h1F;
            16'd32667: data <= 8'h00;
            16'd32668: data <= 8'h1F;
            16'd32669: data <= 8'h00;
            16'd32670: data <= 8'h1F;
            16'd32671: data <= 8'h00;
            16'd32672: data <= 8'h1F;
            16'd32673: data <= 8'h00;
            16'd32674: data <= 8'h1F;
            16'd32675: data <= 8'h00;
            16'd32676: data <= 8'h1F;
            16'd32677: data <= 8'h00;
            16'd32678: data <= 8'h1F;
            16'd32679: data <= 8'h00;
            16'd32680: data <= 8'hFF;
            16'd32681: data <= 8'hFF;
            16'd32682: data <= 8'h1F;
            16'd32683: data <= 8'h00;
            16'd32684: data <= 8'h1F;
            16'd32685: data <= 8'h00;
            16'd32686: data <= 8'h1F;
            16'd32687: data <= 8'h00;
            16'd32688: data <= 8'h1F;
            16'd32689: data <= 8'h00;
            16'd32690: data <= 8'h1F;
            16'd32691: data <= 8'h00;
            16'd32692: data <= 8'h1F;
            16'd32693: data <= 8'h00;
            16'd32694: data <= 8'h1F;
            16'd32695: data <= 8'h00;
            16'd32696: data <= 8'h1F;
            16'd32697: data <= 8'h00;
            16'd32698: data <= 8'h1F;
            16'd32699: data <= 8'h00;
            16'd32700: data <= 8'h1F;
            16'd32701: data <= 8'h00;
            16'd32702: data <= 8'h1F;
            16'd32703: data <= 8'h00;
            16'd32704: data <= 8'h1F;
            16'd32705: data <= 8'h00;
            16'd32706: data <= 8'h1F;
            16'd32707: data <= 8'h00;
            16'd32708: data <= 8'h1F;
            16'd32709: data <= 8'h00;
            16'd32710: data <= 8'h1F;
            16'd32711: data <= 8'h00;
            16'd32712: data <= 8'h1F;
            16'd32713: data <= 8'h00;
            16'd32714: data <= 8'h1F;
            16'd32715: data <= 8'h00;
            16'd32716: data <= 8'h1F;
            16'd32717: data <= 8'h00;
            16'd32718: data <= 8'h1F;
            16'd32719: data <= 8'h00;
            16'd32720: data <= 8'hFF;
            16'd32721: data <= 8'hFF;
            16'd32722: data <= 8'h1F;
            16'd32723: data <= 8'h00;
            16'd32724: data <= 8'h1F;
            16'd32725: data <= 8'h00;
            16'd32726: data <= 8'h1F;
            16'd32727: data <= 8'h00;
            16'd32728: data <= 8'h1F;
            16'd32729: data <= 8'h00;
            16'd32730: data <= 8'h1F;
            16'd32731: data <= 8'h00;
            16'd32732: data <= 8'h1F;
            16'd32733: data <= 8'h00;
            16'd32734: data <= 8'h1F;
            16'd32735: data <= 8'h00;
            16'd32736: data <= 8'h1F;
            16'd32737: data <= 8'h00;
            16'd32738: data <= 8'h1F;
            16'd32739: data <= 8'h00;
            16'd32740: data <= 8'h1F;
            16'd32741: data <= 8'h00;
            16'd32742: data <= 8'h1F;
            16'd32743: data <= 8'h00;
            16'd32744: data <= 8'h1F;
            16'd32745: data <= 8'h00;
            16'd32746: data <= 8'h1F;
            16'd32747: data <= 8'h00;
            16'd32748: data <= 8'h1F;
            16'd32749: data <= 8'h00;
            16'd32750: data <= 8'h1F;
            16'd32751: data <= 8'h00;
            16'd32752: data <= 8'h1F;
            16'd32753: data <= 8'h00;
            16'd32754: data <= 8'h1F;
            16'd32755: data <= 8'h00;
            16'd32756: data <= 8'h1F;
            16'd32757: data <= 8'h00;
            16'd32758: data <= 8'h1F;
            16'd32759: data <= 8'h00;
            16'd32760: data <= 8'hFF;
            16'd32761: data <= 8'hFF;
            16'd32762: data <= 8'h1F;
            16'd32763: data <= 8'h00;
            16'd32764: data <= 8'h1F;
            16'd32765: data <= 8'h00;
            16'd32766: data <= 8'h1F;
            16'd32767: data <= 8'h00;
            16'd32768: data <= 8'h1F;
            16'd32769: data <= 8'h00;
            16'd32770: data <= 8'h1F;
            16'd32771: data <= 8'h00;
            16'd32772: data <= 8'h1F;
            16'd32773: data <= 8'h00;
            16'd32774: data <= 8'h1F;
            16'd32775: data <= 8'h00;
            16'd32776: data <= 8'h1F;
            16'd32777: data <= 8'h00;
            16'd32778: data <= 8'h1F;
            16'd32779: data <= 8'h00;
            16'd32780: data <= 8'h1F;
            16'd32781: data <= 8'h00;
            16'd32782: data <= 8'h1F;
            16'd32783: data <= 8'h00;
            16'd32784: data <= 8'h1F;
            16'd32785: data <= 8'h00;
            16'd32786: data <= 8'h1F;
            16'd32787: data <= 8'h00;
            16'd32788: data <= 8'h1F;
            16'd32789: data <= 8'h00;
            16'd32790: data <= 8'h1F;
            16'd32791: data <= 8'h00;
            16'd32792: data <= 8'h1F;
            16'd32793: data <= 8'h00;
            16'd32794: data <= 8'h1F;
            16'd32795: data <= 8'h00;
            16'd32796: data <= 8'h1F;
            16'd32797: data <= 8'h00;
            16'd32798: data <= 8'h1F;
            16'd32799: data <= 8'h00;
            16'd32800: data <= 8'hFF;
            16'd32801: data <= 8'hFF;
            16'd32802: data <= 8'h1F;
            16'd32803: data <= 8'h00;
            16'd32804: data <= 8'h1F;
            16'd32805: data <= 8'h00;
            16'd32806: data <= 8'h1F;
            16'd32807: data <= 8'h00;
            16'd32808: data <= 8'h1F;
            16'd32809: data <= 8'h00;
            16'd32810: data <= 8'h1F;
            16'd32811: data <= 8'h00;
            16'd32812: data <= 8'h1F;
            16'd32813: data <= 8'h00;
            16'd32814: data <= 8'h1F;
            16'd32815: data <= 8'h00;
            16'd32816: data <= 8'h1F;
            16'd32817: data <= 8'h00;
            16'd32818: data <= 8'h1F;
            16'd32819: data <= 8'h00;
            16'd32820: data <= 8'h1F;
            16'd32821: data <= 8'h00;
            16'd32822: data <= 8'h1F;
            16'd32823: data <= 8'h00;
            16'd32824: data <= 8'h1F;
            16'd32825: data <= 8'h00;
            16'd32826: data <= 8'h1F;
            16'd32827: data <= 8'h00;
            16'd32828: data <= 8'h1F;
            16'd32829: data <= 8'h00;
            16'd32830: data <= 8'h1F;
            16'd32831: data <= 8'h00;
            16'd32832: data <= 8'h1F;
            16'd32833: data <= 8'h00;
            16'd32834: data <= 8'h1F;
            16'd32835: data <= 8'h00;
            16'd32836: data <= 8'h1F;
            16'd32837: data <= 8'h00;
            16'd32838: data <= 8'h1F;
            16'd32839: data <= 8'h00;
            16'd32840: data <= 8'hFF;
            16'd32841: data <= 8'hFF;
            16'd32842: data <= 8'h1F;
            16'd32843: data <= 8'h00;
            16'd32844: data <= 8'h1F;
            16'd32845: data <= 8'h00;
            16'd32846: data <= 8'h1F;
            16'd32847: data <= 8'h00;
            16'd32848: data <= 8'h1F;
            16'd32849: data <= 8'h00;
            16'd32850: data <= 8'h1F;
            16'd32851: data <= 8'h00;
            16'd32852: data <= 8'h1F;
            16'd32853: data <= 8'h00;
            16'd32854: data <= 8'h1F;
            16'd32855: data <= 8'h00;
            16'd32856: data <= 8'h1F;
            16'd32857: data <= 8'h00;
            16'd32858: data <= 8'h1F;
            16'd32859: data <= 8'h00;
            16'd32860: data <= 8'h1F;
            16'd32861: data <= 8'h00;
            16'd32862: data <= 8'h1F;
            16'd32863: data <= 8'h00;
            16'd32864: data <= 8'h1F;
            16'd32865: data <= 8'h00;
            16'd32866: data <= 8'h1F;
            16'd32867: data <= 8'h00;
            16'd32868: data <= 8'h1F;
            16'd32869: data <= 8'h00;
            16'd32870: data <= 8'h1F;
            16'd32871: data <= 8'h00;
            16'd32872: data <= 8'h1F;
            16'd32873: data <= 8'h00;
            16'd32874: data <= 8'h1F;
            16'd32875: data <= 8'h00;
            16'd32876: data <= 8'h1F;
            16'd32877: data <= 8'h00;
            16'd32878: data <= 8'h1F;
            16'd32879: data <= 8'h00;
            16'd32880: data <= 8'hFF;
            16'd32881: data <= 8'hFF;
            16'd32882: data <= 8'h1F;
            16'd32883: data <= 8'h00;
            16'd32884: data <= 8'h1F;
            16'd32885: data <= 8'h00;
            16'd32886: data <= 8'h1F;
            16'd32887: data <= 8'h00;
            16'd32888: data <= 8'h1F;
            16'd32889: data <= 8'h00;
            16'd32890: data <= 8'h1F;
            16'd32891: data <= 8'h00;
            16'd32892: data <= 8'h1F;
            16'd32893: data <= 8'h00;
            16'd32894: data <= 8'h1F;
            16'd32895: data <= 8'h00;
            16'd32896: data <= 8'h1F;
            16'd32897: data <= 8'h00;
            16'd32898: data <= 8'h1F;
            16'd32899: data <= 8'h00;
            16'd32900: data <= 8'h1F;
            16'd32901: data <= 8'h00;
            16'd32902: data <= 8'h1F;
            16'd32903: data <= 8'h00;
            16'd32904: data <= 8'h1F;
            16'd32905: data <= 8'h00;
            16'd32906: data <= 8'h1F;
            16'd32907: data <= 8'h00;
            16'd32908: data <= 8'h1F;
            16'd32909: data <= 8'h00;
            16'd32910: data <= 8'h1F;
            16'd32911: data <= 8'h00;
            16'd32912: data <= 8'h1F;
            16'd32913: data <= 8'h00;
            16'd32914: data <= 8'h1F;
            16'd32915: data <= 8'h00;
            16'd32916: data <= 8'h1F;
            16'd32917: data <= 8'h00;
            16'd32918: data <= 8'h1F;
            16'd32919: data <= 8'h00;
            16'd32920: data <= 8'hFF;
            16'd32921: data <= 8'hFF;
            16'd32922: data <= 8'h1F;
            16'd32923: data <= 8'h00;
            16'd32924: data <= 8'h1F;
            16'd32925: data <= 8'h00;
            16'd32926: data <= 8'h1F;
            16'd32927: data <= 8'h00;
            16'd32928: data <= 8'h1F;
            16'd32929: data <= 8'h00;
            16'd32930: data <= 8'h1F;
            16'd32931: data <= 8'h00;
            16'd32932: data <= 8'h1F;
            16'd32933: data <= 8'h00;
            16'd32934: data <= 8'h1F;
            16'd32935: data <= 8'h00;
            16'd32936: data <= 8'h1F;
            16'd32937: data <= 8'h00;
            16'd32938: data <= 8'h1F;
            16'd32939: data <= 8'h00;
            16'd32940: data <= 8'h1F;
            16'd32941: data <= 8'h00;
            16'd32942: data <= 8'h1F;
            16'd32943: data <= 8'h00;
            16'd32944: data <= 8'h1F;
            16'd32945: data <= 8'h00;
            16'd32946: data <= 8'h1F;
            16'd32947: data <= 8'h00;
            16'd32948: data <= 8'h1F;
            16'd32949: data <= 8'h00;
            16'd32950: data <= 8'h1F;
            16'd32951: data <= 8'h00;
            16'd32952: data <= 8'h1F;
            16'd32953: data <= 8'h00;
            16'd32954: data <= 8'h1F;
            16'd32955: data <= 8'h00;
            16'd32956: data <= 8'h1F;
            16'd32957: data <= 8'h00;
            16'd32958: data <= 8'h1F;
            16'd32959: data <= 8'h00;
            16'd32960: data <= 8'hFF;
            16'd32961: data <= 8'hFF;
            16'd32962: data <= 8'h1F;
            16'd32963: data <= 8'h00;
            16'd32964: data <= 8'h1F;
            16'd32965: data <= 8'h00;
            16'd32966: data <= 8'h1F;
            16'd32967: data <= 8'h00;
            16'd32968: data <= 8'h1F;
            16'd32969: data <= 8'h00;
            16'd32970: data <= 8'h1F;
            16'd32971: data <= 8'h00;
            16'd32972: data <= 8'h1F;
            16'd32973: data <= 8'h00;
            16'd32974: data <= 8'h1F;
            16'd32975: data <= 8'h00;
            16'd32976: data <= 8'h1F;
            16'd32977: data <= 8'h00;
            16'd32978: data <= 8'h1F;
            16'd32979: data <= 8'h00;
            16'd32980: data <= 8'h1F;
            16'd32981: data <= 8'h00;
            16'd32982: data <= 8'h1F;
            16'd32983: data <= 8'h00;
            16'd32984: data <= 8'h1F;
            16'd32985: data <= 8'h00;
            16'd32986: data <= 8'h1F;
            16'd32987: data <= 8'h00;
            16'd32988: data <= 8'h1F;
            16'd32989: data <= 8'h00;
            16'd32990: data <= 8'h1F;
            16'd32991: data <= 8'h00;
            16'd32992: data <= 8'h1F;
            16'd32993: data <= 8'h00;
            16'd32994: data <= 8'h1F;
            16'd32995: data <= 8'h00;
            16'd32996: data <= 8'h1F;
            16'd32997: data <= 8'h00;
            16'd32998: data <= 8'h1F;
            16'd32999: data <= 8'h00;
            16'd33000: data <= 8'hFF;
            16'd33001: data <= 8'hFF;
            16'd33002: data <= 8'h1F;
            16'd33003: data <= 8'h00;
            16'd33004: data <= 8'h1F;
            16'd33005: data <= 8'h00;
            16'd33006: data <= 8'h1F;
            16'd33007: data <= 8'h00;
            16'd33008: data <= 8'h1F;
            16'd33009: data <= 8'h00;
            16'd33010: data <= 8'h1F;
            16'd33011: data <= 8'h00;
            16'd33012: data <= 8'h1F;
            16'd33013: data <= 8'h00;
            16'd33014: data <= 8'h1F;
            16'd33015: data <= 8'h00;
            16'd33016: data <= 8'h1F;
            16'd33017: data <= 8'h00;
            16'd33018: data <= 8'h1F;
            16'd33019: data <= 8'h00;
            16'd33020: data <= 8'h1F;
            16'd33021: data <= 8'h00;
            16'd33022: data <= 8'h1F;
            16'd33023: data <= 8'h00;
            16'd33024: data <= 8'h1F;
            16'd33025: data <= 8'h00;
            16'd33026: data <= 8'h1F;
            16'd33027: data <= 8'h00;
            16'd33028: data <= 8'h1F;
            16'd33029: data <= 8'h00;
            16'd33030: data <= 8'h1F;
            16'd33031: data <= 8'h00;
            16'd33032: data <= 8'h1F;
            16'd33033: data <= 8'h00;
            16'd33034: data <= 8'h1F;
            16'd33035: data <= 8'h00;
            16'd33036: data <= 8'h1F;
            16'd33037: data <= 8'h00;
            16'd33038: data <= 8'h1F;
            16'd33039: data <= 8'h00;
            16'd33040: data <= 8'hFF;
            16'd33041: data <= 8'hFF;
            16'd33042: data <= 8'h1F;
            16'd33043: data <= 8'h00;
            16'd33044: data <= 8'h1F;
            16'd33045: data <= 8'h00;
            16'd33046: data <= 8'h1F;
            16'd33047: data <= 8'h00;
            16'd33048: data <= 8'h1F;
            16'd33049: data <= 8'h00;
            16'd33050: data <= 8'h1F;
            16'd33051: data <= 8'h00;
            16'd33052: data <= 8'h1F;
            16'd33053: data <= 8'h00;
            16'd33054: data <= 8'h1F;
            16'd33055: data <= 8'h00;
            16'd33056: data <= 8'h1F;
            16'd33057: data <= 8'h00;
            16'd33058: data <= 8'h1F;
            16'd33059: data <= 8'h00;
            16'd33060: data <= 8'h1F;
            16'd33061: data <= 8'h00;
            16'd33062: data <= 8'h1F;
            16'd33063: data <= 8'h00;
            16'd33064: data <= 8'h1F;
            16'd33065: data <= 8'h00;
            16'd33066: data <= 8'h1F;
            16'd33067: data <= 8'h00;
            16'd33068: data <= 8'h1F;
            16'd33069: data <= 8'h00;
            16'd33070: data <= 8'h1F;
            16'd33071: data <= 8'h00;
            16'd33072: data <= 8'h1F;
            16'd33073: data <= 8'h00;
            16'd33074: data <= 8'h1F;
            16'd33075: data <= 8'h00;
            16'd33076: data <= 8'h1F;
            16'd33077: data <= 8'h00;
            16'd33078: data <= 8'h1F;
            16'd33079: data <= 8'h00;
            16'd33080: data <= 8'hFF;
            16'd33081: data <= 8'hFF;
            16'd33082: data <= 8'h1F;
            16'd33083: data <= 8'h00;
            16'd33084: data <= 8'h1F;
            16'd33085: data <= 8'h00;
            16'd33086: data <= 8'h1F;
            16'd33087: data <= 8'h00;
            16'd33088: data <= 8'h1F;
            16'd33089: data <= 8'h00;
            16'd33090: data <= 8'h1F;
            16'd33091: data <= 8'h00;
            16'd33092: data <= 8'h1F;
            16'd33093: data <= 8'h00;
            16'd33094: data <= 8'h1F;
            16'd33095: data <= 8'h00;
            16'd33096: data <= 8'h1F;
            16'd33097: data <= 8'h00;
            16'd33098: data <= 8'h1F;
            16'd33099: data <= 8'h00;
            16'd33100: data <= 8'h1F;
            16'd33101: data <= 8'h00;
            16'd33102: data <= 8'h1F;
            16'd33103: data <= 8'h00;
            16'd33104: data <= 8'h1F;
            16'd33105: data <= 8'h00;
            16'd33106: data <= 8'h1F;
            16'd33107: data <= 8'h00;
            16'd33108: data <= 8'h1F;
            16'd33109: data <= 8'h00;
            16'd33110: data <= 8'h1F;
            16'd33111: data <= 8'h00;
            16'd33112: data <= 8'h1F;
            16'd33113: data <= 8'h00;
            16'd33114: data <= 8'h1F;
            16'd33115: data <= 8'h00;
            16'd33116: data <= 8'h1F;
            16'd33117: data <= 8'h00;
            16'd33118: data <= 8'h1F;
            16'd33119: data <= 8'h00;
            16'd33120: data <= 8'hFF;
            16'd33121: data <= 8'hFF;
            16'd33122: data <= 8'h1F;
            16'd33123: data <= 8'h00;
            16'd33124: data <= 8'h1F;
            16'd33125: data <= 8'h00;
            16'd33126: data <= 8'h1F;
            16'd33127: data <= 8'h00;
            16'd33128: data <= 8'h1F;
            16'd33129: data <= 8'h00;
            16'd33130: data <= 8'h1F;
            16'd33131: data <= 8'h00;
            16'd33132: data <= 8'h1F;
            16'd33133: data <= 8'h00;
            16'd33134: data <= 8'h1F;
            16'd33135: data <= 8'h00;
            16'd33136: data <= 8'h1F;
            16'd33137: data <= 8'h00;
            16'd33138: data <= 8'h1F;
            16'd33139: data <= 8'h00;
            16'd33140: data <= 8'h1F;
            16'd33141: data <= 8'h00;
            16'd33142: data <= 8'h1F;
            16'd33143: data <= 8'h00;
            16'd33144: data <= 8'h1F;
            16'd33145: data <= 8'h00;
            16'd33146: data <= 8'h1F;
            16'd33147: data <= 8'h00;
            16'd33148: data <= 8'h1F;
            16'd33149: data <= 8'h00;
            16'd33150: data <= 8'h1F;
            16'd33151: data <= 8'h00;
            16'd33152: data <= 8'h1F;
            16'd33153: data <= 8'h00;
            16'd33154: data <= 8'h1F;
            16'd33155: data <= 8'h00;
            16'd33156: data <= 8'h1F;
            16'd33157: data <= 8'h00;
            16'd33158: data <= 8'h1F;
            16'd33159: data <= 8'h00;
            16'd33160: data <= 8'hFF;
            16'd33161: data <= 8'hFF;
            16'd33162: data <= 8'h1F;
            16'd33163: data <= 8'h00;
            16'd33164: data <= 8'h1F;
            16'd33165: data <= 8'h00;
            16'd33166: data <= 8'h1F;
            16'd33167: data <= 8'h00;
            16'd33168: data <= 8'h1F;
            16'd33169: data <= 8'h00;
            16'd33170: data <= 8'h1F;
            16'd33171: data <= 8'h00;
            16'd33172: data <= 8'h1F;
            16'd33173: data <= 8'h00;
            16'd33174: data <= 8'h1F;
            16'd33175: data <= 8'h00;
            16'd33176: data <= 8'h1F;
            16'd33177: data <= 8'h00;
            16'd33178: data <= 8'h1F;
            16'd33179: data <= 8'h00;
            16'd33180: data <= 8'h1F;
            16'd33181: data <= 8'h00;
            16'd33182: data <= 8'h1F;
            16'd33183: data <= 8'h00;
            16'd33184: data <= 8'h1F;
            16'd33185: data <= 8'h00;
            16'd33186: data <= 8'h1F;
            16'd33187: data <= 8'h00;
            16'd33188: data <= 8'h1F;
            16'd33189: data <= 8'h00;
            16'd33190: data <= 8'h1F;
            16'd33191: data <= 8'h00;
            16'd33192: data <= 8'h1F;
            16'd33193: data <= 8'h00;
            16'd33194: data <= 8'h1F;
            16'd33195: data <= 8'h00;
            16'd33196: data <= 8'h1F;
            16'd33197: data <= 8'h00;
            16'd33198: data <= 8'h1F;
            16'd33199: data <= 8'h00;
            16'd33200: data <= 8'hFF;
            16'd33201: data <= 8'hFF;
            16'd33202: data <= 8'h1F;
            16'd33203: data <= 8'h00;
            16'd33204: data <= 8'h1F;
            16'd33205: data <= 8'h00;
            16'd33206: data <= 8'h1F;
            16'd33207: data <= 8'h00;
            16'd33208: data <= 8'h1F;
            16'd33209: data <= 8'h00;
            16'd33210: data <= 8'h1F;
            16'd33211: data <= 8'h00;
            16'd33212: data <= 8'h1F;
            16'd33213: data <= 8'h00;
            16'd33214: data <= 8'h1F;
            16'd33215: data <= 8'h00;
            16'd33216: data <= 8'h1F;
            16'd33217: data <= 8'h00;
            16'd33218: data <= 8'h1F;
            16'd33219: data <= 8'h00;
            16'd33220: data <= 8'h1F;
            16'd33221: data <= 8'h00;
            16'd33222: data <= 8'h1F;
            16'd33223: data <= 8'h00;
            16'd33224: data <= 8'h1F;
            16'd33225: data <= 8'h00;
            16'd33226: data <= 8'h1F;
            16'd33227: data <= 8'h00;
            16'd33228: data <= 8'h1F;
            16'd33229: data <= 8'h00;
            16'd33230: data <= 8'h1F;
            16'd33231: data <= 8'h00;
            16'd33232: data <= 8'h1F;
            16'd33233: data <= 8'h00;
            16'd33234: data <= 8'h1F;
            16'd33235: data <= 8'h00;
            16'd33236: data <= 8'h1F;
            16'd33237: data <= 8'h00;
            16'd33238: data <= 8'h1F;
            16'd33239: data <= 8'h00;
            16'd33240: data <= 8'hFF;
            16'd33241: data <= 8'hFF;
            16'd33242: data <= 8'h1F;
            16'd33243: data <= 8'h00;
            16'd33244: data <= 8'h1F;
            16'd33245: data <= 8'h00;
            16'd33246: data <= 8'h1F;
            16'd33247: data <= 8'h00;
            16'd33248: data <= 8'h1F;
            16'd33249: data <= 8'h00;
            16'd33250: data <= 8'h1F;
            16'd33251: data <= 8'h00;
            16'd33252: data <= 8'h1F;
            16'd33253: data <= 8'h00;
            16'd33254: data <= 8'h1F;
            16'd33255: data <= 8'h00;
            16'd33256: data <= 8'h1F;
            16'd33257: data <= 8'h00;
            16'd33258: data <= 8'h1F;
            16'd33259: data <= 8'h00;
            16'd33260: data <= 8'h1F;
            16'd33261: data <= 8'h00;
            16'd33262: data <= 8'h1F;
            16'd33263: data <= 8'h00;
            16'd33264: data <= 8'h1F;
            16'd33265: data <= 8'h00;
            16'd33266: data <= 8'h1F;
            16'd33267: data <= 8'h00;
            16'd33268: data <= 8'h1F;
            16'd33269: data <= 8'h00;
            16'd33270: data <= 8'h1F;
            16'd33271: data <= 8'h00;
            16'd33272: data <= 8'h1F;
            16'd33273: data <= 8'h00;
            16'd33274: data <= 8'h1F;
            16'd33275: data <= 8'h00;
            16'd33276: data <= 8'h1F;
            16'd33277: data <= 8'h00;
            16'd33278: data <= 8'h1F;
            16'd33279: data <= 8'h00;
            16'd33280: data <= 8'hFF;
            16'd33281: data <= 8'hFF;
            16'd33282: data <= 8'h1F;
            16'd33283: data <= 8'h00;
            16'd33284: data <= 8'h1F;
            16'd33285: data <= 8'h00;
            16'd33286: data <= 8'h1F;
            16'd33287: data <= 8'h00;
            16'd33288: data <= 8'h1F;
            16'd33289: data <= 8'h00;
            16'd33290: data <= 8'h1F;
            16'd33291: data <= 8'h00;
            16'd33292: data <= 8'h1F;
            16'd33293: data <= 8'h00;
            16'd33294: data <= 8'h1F;
            16'd33295: data <= 8'h00;
            16'd33296: data <= 8'h1F;
            16'd33297: data <= 8'h00;
            16'd33298: data <= 8'h1F;
            16'd33299: data <= 8'h00;
            16'd33300: data <= 8'h1F;
            16'd33301: data <= 8'h00;
            16'd33302: data <= 8'h1F;
            16'd33303: data <= 8'h00;
            16'd33304: data <= 8'h1F;
            16'd33305: data <= 8'h00;
            16'd33306: data <= 8'h1F;
            16'd33307: data <= 8'h00;
            16'd33308: data <= 8'h1F;
            16'd33309: data <= 8'h00;
            16'd33310: data <= 8'h1F;
            16'd33311: data <= 8'h00;
            16'd33312: data <= 8'h1F;
            16'd33313: data <= 8'h00;
            16'd33314: data <= 8'h1F;
            16'd33315: data <= 8'h00;
            16'd33316: data <= 8'h1F;
            16'd33317: data <= 8'h00;
            16'd33318: data <= 8'h1F;
            16'd33319: data <= 8'h00;
            16'd33320: data <= 8'hFF;
            16'd33321: data <= 8'hFF;
            16'd33322: data <= 8'h1F;
            16'd33323: data <= 8'h00;
            16'd33324: data <= 8'h1F;
            16'd33325: data <= 8'h00;
            16'd33326: data <= 8'h1F;
            16'd33327: data <= 8'h00;
            16'd33328: data <= 8'h1F;
            16'd33329: data <= 8'h00;
            16'd33330: data <= 8'h1F;
            16'd33331: data <= 8'h00;
            16'd33332: data <= 8'h1F;
            16'd33333: data <= 8'h00;
            16'd33334: data <= 8'h1F;
            16'd33335: data <= 8'h00;
            16'd33336: data <= 8'h1F;
            16'd33337: data <= 8'h00;
            16'd33338: data <= 8'h1F;
            16'd33339: data <= 8'h00;
            16'd33340: data <= 8'h1F;
            16'd33341: data <= 8'h00;
            16'd33342: data <= 8'h1F;
            16'd33343: data <= 8'h00;
            16'd33344: data <= 8'h1F;
            16'd33345: data <= 8'h00;
            16'd33346: data <= 8'h1F;
            16'd33347: data <= 8'h00;
            16'd33348: data <= 8'h1F;
            16'd33349: data <= 8'h00;
            16'd33350: data <= 8'h1F;
            16'd33351: data <= 8'h00;
            16'd33352: data <= 8'h1F;
            16'd33353: data <= 8'h00;
            16'd33354: data <= 8'h1F;
            16'd33355: data <= 8'h00;
            16'd33356: data <= 8'h1F;
            16'd33357: data <= 8'h00;
            16'd33358: data <= 8'h1F;
            16'd33359: data <= 8'h00;
            16'd33360: data <= 8'hFF;
            16'd33361: data <= 8'hFF;
            16'd33362: data <= 8'h1F;
            16'd33363: data <= 8'h00;
            16'd33364: data <= 8'h1F;
            16'd33365: data <= 8'h00;
            16'd33366: data <= 8'h1F;
            16'd33367: data <= 8'h00;
            16'd33368: data <= 8'h1F;
            16'd33369: data <= 8'h00;
            16'd33370: data <= 8'h1F;
            16'd33371: data <= 8'h00;
            16'd33372: data <= 8'h1F;
            16'd33373: data <= 8'h00;
            16'd33374: data <= 8'h1F;
            16'd33375: data <= 8'h00;
            16'd33376: data <= 8'h1F;
            16'd33377: data <= 8'h00;
            16'd33378: data <= 8'h1F;
            16'd33379: data <= 8'h00;
            16'd33380: data <= 8'h1F;
            16'd33381: data <= 8'h00;
            16'd33382: data <= 8'h1F;
            16'd33383: data <= 8'h00;
            16'd33384: data <= 8'h1F;
            16'd33385: data <= 8'h00;
            16'd33386: data <= 8'h1F;
            16'd33387: data <= 8'h00;
            16'd33388: data <= 8'h1F;
            16'd33389: data <= 8'h00;
            16'd33390: data <= 8'h1F;
            16'd33391: data <= 8'h00;
            16'd33392: data <= 8'h1F;
            16'd33393: data <= 8'h00;
            16'd33394: data <= 8'h1F;
            16'd33395: data <= 8'h00;
            16'd33396: data <= 8'h1F;
            16'd33397: data <= 8'h00;
            16'd33398: data <= 8'h1F;
            16'd33399: data <= 8'h00;
            16'd33400: data <= 8'hFF;
            16'd33401: data <= 8'hFF;
            16'd33402: data <= 8'h1F;
            16'd33403: data <= 8'h00;
            16'd33404: data <= 8'h1F;
            16'd33405: data <= 8'h00;
            16'd33406: data <= 8'h1F;
            16'd33407: data <= 8'h00;
            16'd33408: data <= 8'h1F;
            16'd33409: data <= 8'h00;
            16'd33410: data <= 8'h1F;
            16'd33411: data <= 8'h00;
            16'd33412: data <= 8'h1F;
            16'd33413: data <= 8'h00;
            16'd33414: data <= 8'h1F;
            16'd33415: data <= 8'h00;
            16'd33416: data <= 8'h1F;
            16'd33417: data <= 8'h00;
            16'd33418: data <= 8'h1F;
            16'd33419: data <= 8'h00;
            16'd33420: data <= 8'h1F;
            16'd33421: data <= 8'h00;
            16'd33422: data <= 8'h1F;
            16'd33423: data <= 8'h00;
            16'd33424: data <= 8'h1F;
            16'd33425: data <= 8'h00;
            16'd33426: data <= 8'h1F;
            16'd33427: data <= 8'h00;
            16'd33428: data <= 8'h1F;
            16'd33429: data <= 8'h00;
            16'd33430: data <= 8'h1F;
            16'd33431: data <= 8'h00;
            16'd33432: data <= 8'h1F;
            16'd33433: data <= 8'h00;
            16'd33434: data <= 8'h1F;
            16'd33435: data <= 8'h00;
            16'd33436: data <= 8'h1F;
            16'd33437: data <= 8'h00;
            16'd33438: data <= 8'h1F;
            16'd33439: data <= 8'h00;
            16'd33440: data <= 8'hFF;
            16'd33441: data <= 8'hFF;
            16'd33442: data <= 8'h1F;
            16'd33443: data <= 8'h00;
            16'd33444: data <= 8'h1F;
            16'd33445: data <= 8'h00;
            16'd33446: data <= 8'h1F;
            16'd33447: data <= 8'h00;
            16'd33448: data <= 8'h1F;
            16'd33449: data <= 8'h00;
            16'd33450: data <= 8'h1F;
            16'd33451: data <= 8'h00;
            16'd33452: data <= 8'h1F;
            16'd33453: data <= 8'h00;
            16'd33454: data <= 8'h1F;
            16'd33455: data <= 8'h00;
            16'd33456: data <= 8'h1F;
            16'd33457: data <= 8'h00;
            16'd33458: data <= 8'h1F;
            16'd33459: data <= 8'h00;
            16'd33460: data <= 8'h1F;
            16'd33461: data <= 8'h00;
            16'd33462: data <= 8'h1F;
            16'd33463: data <= 8'h00;
            16'd33464: data <= 8'h1F;
            16'd33465: data <= 8'h00;
            16'd33466: data <= 8'h1F;
            16'd33467: data <= 8'h00;
            16'd33468: data <= 8'h1F;
            16'd33469: data <= 8'h00;
            16'd33470: data <= 8'h1F;
            16'd33471: data <= 8'h00;
            16'd33472: data <= 8'h1F;
            16'd33473: data <= 8'h00;
            16'd33474: data <= 8'h1F;
            16'd33475: data <= 8'h00;
            16'd33476: data <= 8'h1F;
            16'd33477: data <= 8'h00;
            16'd33478: data <= 8'h1F;
            16'd33479: data <= 8'h00;
            16'd33480: data <= 8'hFF;
            16'd33481: data <= 8'hFF;
            16'd33482: data <= 8'h1F;
            16'd33483: data <= 8'h00;
            16'd33484: data <= 8'h1F;
            16'd33485: data <= 8'h00;
            16'd33486: data <= 8'h1F;
            16'd33487: data <= 8'h00;
            16'd33488: data <= 8'h1F;
            16'd33489: data <= 8'h00;
            16'd33490: data <= 8'h1F;
            16'd33491: data <= 8'h00;
            16'd33492: data <= 8'h1F;
            16'd33493: data <= 8'h00;
            16'd33494: data <= 8'h1F;
            16'd33495: data <= 8'h00;
            16'd33496: data <= 8'h1F;
            16'd33497: data <= 8'h00;
            16'd33498: data <= 8'h1F;
            16'd33499: data <= 8'h00;
            16'd33500: data <= 8'h1F;
            16'd33501: data <= 8'h00;
            16'd33502: data <= 8'h1F;
            16'd33503: data <= 8'h00;
            16'd33504: data <= 8'h1F;
            16'd33505: data <= 8'h00;
            16'd33506: data <= 8'h1F;
            16'd33507: data <= 8'h00;
            16'd33508: data <= 8'h1F;
            16'd33509: data <= 8'h00;
            16'd33510: data <= 8'h1F;
            16'd33511: data <= 8'h00;
            16'd33512: data <= 8'h1F;
            16'd33513: data <= 8'h00;
            16'd33514: data <= 8'h1F;
            16'd33515: data <= 8'h00;
            16'd33516: data <= 8'h1F;
            16'd33517: data <= 8'h00;
            16'd33518: data <= 8'h1F;
            16'd33519: data <= 8'h00;
            16'd33520: data <= 8'hFF;
            16'd33521: data <= 8'hFF;
            16'd33522: data <= 8'h1F;
            16'd33523: data <= 8'h00;
            16'd33524: data <= 8'h1F;
            16'd33525: data <= 8'h00;
            16'd33526: data <= 8'h1F;
            16'd33527: data <= 8'h00;
            16'd33528: data <= 8'h1F;
            16'd33529: data <= 8'h00;
            16'd33530: data <= 8'h1F;
            16'd33531: data <= 8'h00;
            16'd33532: data <= 8'h1F;
            16'd33533: data <= 8'h00;
            16'd33534: data <= 8'h1F;
            16'd33535: data <= 8'h00;
            16'd33536: data <= 8'h1F;
            16'd33537: data <= 8'h00;
            16'd33538: data <= 8'h1F;
            16'd33539: data <= 8'h00;
            16'd33540: data <= 8'h1F;
            16'd33541: data <= 8'h00;
            16'd33542: data <= 8'h1F;
            16'd33543: data <= 8'h00;
            16'd33544: data <= 8'h1F;
            16'd33545: data <= 8'h00;
            16'd33546: data <= 8'h1F;
            16'd33547: data <= 8'h00;
            16'd33548: data <= 8'h1F;
            16'd33549: data <= 8'h00;
            16'd33550: data <= 8'h1F;
            16'd33551: data <= 8'h00;
            16'd33552: data <= 8'h1F;
            16'd33553: data <= 8'h00;
            16'd33554: data <= 8'h1F;
            16'd33555: data <= 8'h00;
            16'd33556: data <= 8'h1F;
            16'd33557: data <= 8'h00;
            16'd33558: data <= 8'h1F;
            16'd33559: data <= 8'h00;
            16'd33560: data <= 8'hFF;
            16'd33561: data <= 8'hFF;
            16'd33562: data <= 8'h1F;
            16'd33563: data <= 8'h00;
            16'd33564: data <= 8'h1F;
            16'd33565: data <= 8'h00;
            16'd33566: data <= 8'h1F;
            16'd33567: data <= 8'h00;
            16'd33568: data <= 8'h1F;
            16'd33569: data <= 8'h00;
            16'd33570: data <= 8'h1F;
            16'd33571: data <= 8'h00;
            16'd33572: data <= 8'h1F;
            16'd33573: data <= 8'h00;
            16'd33574: data <= 8'h1F;
            16'd33575: data <= 8'h00;
            16'd33576: data <= 8'h1F;
            16'd33577: data <= 8'h00;
            16'd33578: data <= 8'h1F;
            16'd33579: data <= 8'h00;
            16'd33580: data <= 8'h1F;
            16'd33581: data <= 8'h00;
            16'd33582: data <= 8'h1F;
            16'd33583: data <= 8'h00;
            16'd33584: data <= 8'h1F;
            16'd33585: data <= 8'h00;
            16'd33586: data <= 8'h1F;
            16'd33587: data <= 8'h00;
            16'd33588: data <= 8'h1F;
            16'd33589: data <= 8'h00;
            16'd33590: data <= 8'h1F;
            16'd33591: data <= 8'h00;
            16'd33592: data <= 8'h1F;
            16'd33593: data <= 8'h00;
            16'd33594: data <= 8'h1F;
            16'd33595: data <= 8'h00;
            16'd33596: data <= 8'h1F;
            16'd33597: data <= 8'h00;
            16'd33598: data <= 8'h1F;
            16'd33599: data <= 8'h00;
            16'd33600: data <= 8'hFF;
            16'd33601: data <= 8'hFF;
            16'd33602: data <= 8'hFF;
            16'd33603: data <= 8'hFF;
            16'd33604: data <= 8'hFF;
            16'd33605: data <= 8'hFF;
            16'd33606: data <= 8'hFF;
            16'd33607: data <= 8'hFF;
            16'd33608: data <= 8'hFF;
            16'd33609: data <= 8'hFF;
            16'd33610: data <= 8'hFF;
            16'd33611: data <= 8'hFF;
            16'd33612: data <= 8'hFF;
            16'd33613: data <= 8'hFF;
            16'd33614: data <= 8'hFF;
            16'd33615: data <= 8'hFF;
            16'd33616: data <= 8'hFF;
            16'd33617: data <= 8'hFF;
            16'd33618: data <= 8'hFF;
            16'd33619: data <= 8'hFF;
            16'd33620: data <= 8'hFF;
            16'd33621: data <= 8'hFF;
            16'd33622: data <= 8'hFF;
            16'd33623: data <= 8'hFF;
            16'd33624: data <= 8'hFF;
            16'd33625: data <= 8'hFF;
            16'd33626: data <= 8'hFF;
            16'd33627: data <= 8'hFF;
            16'd33628: data <= 8'hFF;
            16'd33629: data <= 8'hFF;
            16'd33630: data <= 8'hFF;
            16'd33631: data <= 8'hFF;
            16'd33632: data <= 8'hFF;
            16'd33633: data <= 8'hFF;
            16'd33634: data <= 8'hFF;
            16'd33635: data <= 8'hFF;
            16'd33636: data <= 8'hFF;
            16'd33637: data <= 8'hFF;
            16'd33638: data <= 8'hFF;
            16'd33639: data <= 8'hFF;
            16'd33640: data <= 8'hFF;
            16'd33641: data <= 8'hFF;
            16'd33642: data <= 8'hFF;
            16'd33643: data <= 8'hFF;
            16'd33644: data <= 8'hFF;
            16'd33645: data <= 8'hFF;
            16'd33646: data <= 8'hFF;
            16'd33647: data <= 8'hFF;
            16'd33648: data <= 8'hFF;
            16'd33649: data <= 8'hFF;
            16'd33650: data <= 8'hFF;
            16'd33651: data <= 8'hFF;
            16'd33652: data <= 8'hFF;
            16'd33653: data <= 8'hFF;
            16'd33654: data <= 8'hFF;
            16'd33655: data <= 8'hFF;
            16'd33656: data <= 8'hFF;
            16'd33657: data <= 8'hFF;
            16'd33658: data <= 8'hFF;
            16'd33659: data <= 8'hFF;
            16'd33660: data <= 8'hFF;
            16'd33661: data <= 8'hFF;
            16'd33662: data <= 8'hFF;
            16'd33663: data <= 8'hFF;
            16'd33664: data <= 8'hFF;
            16'd33665: data <= 8'hFF;
            16'd33666: data <= 8'hFF;
            16'd33667: data <= 8'hFF;
            16'd33668: data <= 8'hFF;
            16'd33669: data <= 8'hFF;
            16'd33670: data <= 8'hFF;
            16'd33671: data <= 8'hFF;
            16'd33672: data <= 8'hFF;
            16'd33673: data <= 8'hFF;
            16'd33674: data <= 8'hFF;
            16'd33675: data <= 8'hFF;
            16'd33676: data <= 8'hFF;
            16'd33677: data <= 8'hFF;
            16'd33678: data <= 8'hFF;
            16'd33679: data <= 8'hFF;
            16'd33680: data <= 8'hFF;
            16'd33681: data <= 8'hFF;
            16'd33682: data <= 8'hFF;
            16'd33683: data <= 8'hFF;
            16'd33684: data <= 8'hFF;
            16'd33685: data <= 8'hFF;
            16'd33686: data <= 8'hFF;
            16'd33687: data <= 8'hFF;
            16'd33688: data <= 8'hFF;
            16'd33689: data <= 8'hFF;
            16'd33690: data <= 8'hFF;
            16'd33691: data <= 8'hFF;
            16'd33692: data <= 8'hFF;
            16'd33693: data <= 8'hFF;
            16'd33694: data <= 8'hFF;
            16'd33695: data <= 8'hFF;
            16'd33696: data <= 8'hFF;
            16'd33697: data <= 8'hFF;
            16'd33698: data <= 8'hFF;
            16'd33699: data <= 8'hFF;
            16'd33700: data <= 8'hFF;
            16'd33701: data <= 8'hFF;
            16'd33702: data <= 8'hFF;
            16'd33703: data <= 8'hFF;
            16'd33704: data <= 8'hFF;
            16'd33705: data <= 8'hFF;
            16'd33706: data <= 8'hFF;
            16'd33707: data <= 8'hFF;
            16'd33708: data <= 8'hFF;
            16'd33709: data <= 8'hFF;
            16'd33710: data <= 8'hFF;
            16'd33711: data <= 8'hFF;
            16'd33712: data <= 8'hFF;
            16'd33713: data <= 8'hFF;
            16'd33714: data <= 8'hFF;
            16'd33715: data <= 8'hFF;
            16'd33716: data <= 8'hFF;
            16'd33717: data <= 8'hFF;
            16'd33718: data <= 8'hFF;
            16'd33719: data <= 8'hFF;
            16'd33720: data <= 8'hFF;
            16'd33721: data <= 8'hFF;
            16'd33722: data <= 8'hFF;
            16'd33723: data <= 8'hFF;
            16'd33724: data <= 8'hFF;
            16'd33725: data <= 8'hFF;
            16'd33726: data <= 8'hFF;
            16'd33727: data <= 8'hFF;
            16'd33728: data <= 8'hFF;
            16'd33729: data <= 8'hFF;
            16'd33730: data <= 8'hFF;
            16'd33731: data <= 8'hFF;
            16'd33732: data <= 8'hFF;
            16'd33733: data <= 8'hFF;
            16'd33734: data <= 8'hFF;
            16'd33735: data <= 8'hFF;
            16'd33736: data <= 8'hFF;
            16'd33737: data <= 8'hFF;
            16'd33738: data <= 8'hFF;
            16'd33739: data <= 8'hFF;
            16'd33740: data <= 8'hFF;
            16'd33741: data <= 8'hFF;
            16'd33742: data <= 8'hFF;
            16'd33743: data <= 8'hFF;
            16'd33744: data <= 8'hFF;
            16'd33745: data <= 8'hFF;
            16'd33746: data <= 8'hFF;
            16'd33747: data <= 8'hFF;
            16'd33748: data <= 8'hFF;
            16'd33749: data <= 8'hFF;
            16'd33750: data <= 8'hFF;
            16'd33751: data <= 8'hFF;
            16'd33752: data <= 8'hFF;
            16'd33753: data <= 8'hFF;
            16'd33754: data <= 8'hFF;
            16'd33755: data <= 8'hFF;
            16'd33756: data <= 8'hFF;
            16'd33757: data <= 8'hFF;
            16'd33758: data <= 8'hFF;
            16'd33759: data <= 8'hFF;
            16'd33760: data <= 8'hFF;
            16'd33761: data <= 8'hFF;
            16'd33762: data <= 8'hFF;
            16'd33763: data <= 8'hFF;
            16'd33764: data <= 8'hFF;
            16'd33765: data <= 8'hFF;
            16'd33766: data <= 8'hFF;
            16'd33767: data <= 8'hFF;
            16'd33768: data <= 8'hFF;
            16'd33769: data <= 8'hFF;
            16'd33770: data <= 8'hFF;
            16'd33771: data <= 8'hFF;
            16'd33772: data <= 8'hFF;
            16'd33773: data <= 8'hFF;
            16'd33774: data <= 8'hFF;
            16'd33775: data <= 8'hFF;
            16'd33776: data <= 8'hFF;
            16'd33777: data <= 8'hFF;
            16'd33778: data <= 8'hFF;
            16'd33779: data <= 8'hFF;
            16'd33780: data <= 8'hFF;
            16'd33781: data <= 8'hFF;
            16'd33782: data <= 8'hFF;
            16'd33783: data <= 8'hFF;
            16'd33784: data <= 8'hFF;
            16'd33785: data <= 8'hFF;
            16'd33786: data <= 8'hFF;
            16'd33787: data <= 8'hFF;
            16'd33788: data <= 8'hFF;
            16'd33789: data <= 8'hFF;
            16'd33790: data <= 8'hFF;
            16'd33791: data <= 8'hFF;
            16'd33792: data <= 8'hFF;
            16'd33793: data <= 8'hFF;
            16'd33794: data <= 8'hFF;
            16'd33795: data <= 8'hFF;
            16'd33796: data <= 8'hFF;
            16'd33797: data <= 8'hFF;
            16'd33798: data <= 8'hFF;
            16'd33799: data <= 8'hFF;
            16'd33800: data <= 8'hFF;
            16'd33801: data <= 8'hFF;
            16'd33802: data <= 8'hFF;
            16'd33803: data <= 8'hFF;
            16'd33804: data <= 8'hFF;
            16'd33805: data <= 8'hFF;
            16'd33806: data <= 8'hFF;
            16'd33807: data <= 8'hFF;
            16'd33808: data <= 8'hFF;
            16'd33809: data <= 8'hFF;
            16'd33810: data <= 8'hFF;
            16'd33811: data <= 8'hFF;
            16'd33812: data <= 8'hFF;
            16'd33813: data <= 8'hFF;
            16'd33814: data <= 8'hFF;
            16'd33815: data <= 8'hFF;
            16'd33816: data <= 8'hFF;
            16'd33817: data <= 8'hFF;
            16'd33818: data <= 8'hFF;
            16'd33819: data <= 8'hFF;
            16'd33820: data <= 8'hFF;
            16'd33821: data <= 8'hFF;
            16'd33822: data <= 8'hFF;
            16'd33823: data <= 8'hFF;
            16'd33824: data <= 8'hFF;
            16'd33825: data <= 8'hFF;
            16'd33826: data <= 8'hFF;
            16'd33827: data <= 8'hFF;
            16'd33828: data <= 8'hFF;
            16'd33829: data <= 8'hFF;
            16'd33830: data <= 8'hFF;
            16'd33831: data <= 8'hFF;
            16'd33832: data <= 8'hFF;
            16'd33833: data <= 8'hFF;
            16'd33834: data <= 8'hFF;
            16'd33835: data <= 8'hFF;
            16'd33836: data <= 8'hFF;
            16'd33837: data <= 8'hFF;
            16'd33838: data <= 8'hFF;
            16'd33839: data <= 8'hFF;
            16'd33840: data <= 8'hFF;
            16'd33841: data <= 8'hFF;
            16'd33842: data <= 8'h1F;
            16'd33843: data <= 8'h00;
            16'd33844: data <= 8'h1F;
            16'd33845: data <= 8'h00;
            16'd33846: data <= 8'h1F;
            16'd33847: data <= 8'h00;
            16'd33848: data <= 8'h1F;
            16'd33849: data <= 8'h00;
            16'd33850: data <= 8'h1F;
            16'd33851: data <= 8'h00;
            16'd33852: data <= 8'h1F;
            16'd33853: data <= 8'h00;
            16'd33854: data <= 8'h1F;
            16'd33855: data <= 8'h00;
            16'd33856: data <= 8'h1F;
            16'd33857: data <= 8'h00;
            16'd33858: data <= 8'h1F;
            16'd33859: data <= 8'h00;
            16'd33860: data <= 8'h1F;
            16'd33861: data <= 8'h00;
            16'd33862: data <= 8'h1F;
            16'd33863: data <= 8'h00;
            16'd33864: data <= 8'h1F;
            16'd33865: data <= 8'h00;
            16'd33866: data <= 8'h1F;
            16'd33867: data <= 8'h00;
            16'd33868: data <= 8'h1F;
            16'd33869: data <= 8'h00;
            16'd33870: data <= 8'h1F;
            16'd33871: data <= 8'h00;
            16'd33872: data <= 8'h1F;
            16'd33873: data <= 8'h00;
            16'd33874: data <= 8'h1F;
            16'd33875: data <= 8'h00;
            16'd33876: data <= 8'h1F;
            16'd33877: data <= 8'h00;
            16'd33878: data <= 8'h1F;
            16'd33879: data <= 8'h00;
            16'd33880: data <= 8'hFF;
            16'd33881: data <= 8'hFF;
            16'd33882: data <= 8'h1F;
            16'd33883: data <= 8'h00;
            16'd33884: data <= 8'h1F;
            16'd33885: data <= 8'h00;
            16'd33886: data <= 8'h1F;
            16'd33887: data <= 8'h00;
            16'd33888: data <= 8'h1F;
            16'd33889: data <= 8'h00;
            16'd33890: data <= 8'h1F;
            16'd33891: data <= 8'h00;
            16'd33892: data <= 8'h1F;
            16'd33893: data <= 8'h00;
            16'd33894: data <= 8'h1F;
            16'd33895: data <= 8'h00;
            16'd33896: data <= 8'h1F;
            16'd33897: data <= 8'h00;
            16'd33898: data <= 8'h1F;
            16'd33899: data <= 8'h00;
            16'd33900: data <= 8'h1F;
            16'd33901: data <= 8'h00;
            16'd33902: data <= 8'h1F;
            16'd33903: data <= 8'h00;
            16'd33904: data <= 8'h1F;
            16'd33905: data <= 8'h00;
            16'd33906: data <= 8'h1F;
            16'd33907: data <= 8'h00;
            16'd33908: data <= 8'h1F;
            16'd33909: data <= 8'h00;
            16'd33910: data <= 8'h1F;
            16'd33911: data <= 8'h00;
            16'd33912: data <= 8'h1F;
            16'd33913: data <= 8'h00;
            16'd33914: data <= 8'h1F;
            16'd33915: data <= 8'h00;
            16'd33916: data <= 8'h1F;
            16'd33917: data <= 8'h00;
            16'd33918: data <= 8'h1F;
            16'd33919: data <= 8'h00;
            16'd33920: data <= 8'hFF;
            16'd33921: data <= 8'hFF;
            16'd33922: data <= 8'h1F;
            16'd33923: data <= 8'h00;
            16'd33924: data <= 8'h1F;
            16'd33925: data <= 8'h00;
            16'd33926: data <= 8'h1F;
            16'd33927: data <= 8'h00;
            16'd33928: data <= 8'h1F;
            16'd33929: data <= 8'h00;
            16'd33930: data <= 8'h1F;
            16'd33931: data <= 8'h00;
            16'd33932: data <= 8'h1F;
            16'd33933: data <= 8'h00;
            16'd33934: data <= 8'h1F;
            16'd33935: data <= 8'h00;
            16'd33936: data <= 8'h1F;
            16'd33937: data <= 8'h00;
            16'd33938: data <= 8'h1F;
            16'd33939: data <= 8'h00;
            16'd33940: data <= 8'h1F;
            16'd33941: data <= 8'h00;
            16'd33942: data <= 8'h1F;
            16'd33943: data <= 8'h00;
            16'd33944: data <= 8'h1F;
            16'd33945: data <= 8'h00;
            16'd33946: data <= 8'h1F;
            16'd33947: data <= 8'h00;
            16'd33948: data <= 8'h1F;
            16'd33949: data <= 8'h00;
            16'd33950: data <= 8'h1F;
            16'd33951: data <= 8'h00;
            16'd33952: data <= 8'h1F;
            16'd33953: data <= 8'h00;
            16'd33954: data <= 8'h1F;
            16'd33955: data <= 8'h00;
            16'd33956: data <= 8'h1F;
            16'd33957: data <= 8'h00;
            16'd33958: data <= 8'h1F;
            16'd33959: data <= 8'h00;
            16'd33960: data <= 8'hFF;
            16'd33961: data <= 8'hFF;
            16'd33962: data <= 8'h1F;
            16'd33963: data <= 8'h00;
            16'd33964: data <= 8'h1F;
            16'd33965: data <= 8'h00;
            16'd33966: data <= 8'h1F;
            16'd33967: data <= 8'h00;
            16'd33968: data <= 8'h1F;
            16'd33969: data <= 8'h00;
            16'd33970: data <= 8'h1F;
            16'd33971: data <= 8'h00;
            16'd33972: data <= 8'h1F;
            16'd33973: data <= 8'h00;
            16'd33974: data <= 8'h1F;
            16'd33975: data <= 8'h00;
            16'd33976: data <= 8'h1F;
            16'd33977: data <= 8'h00;
            16'd33978: data <= 8'h1F;
            16'd33979: data <= 8'h00;
            16'd33980: data <= 8'h1F;
            16'd33981: data <= 8'h00;
            16'd33982: data <= 8'h1F;
            16'd33983: data <= 8'h00;
            16'd33984: data <= 8'h1F;
            16'd33985: data <= 8'h00;
            16'd33986: data <= 8'h1F;
            16'd33987: data <= 8'h00;
            16'd33988: data <= 8'h1F;
            16'd33989: data <= 8'h00;
            16'd33990: data <= 8'h1F;
            16'd33991: data <= 8'h00;
            16'd33992: data <= 8'h1F;
            16'd33993: data <= 8'h00;
            16'd33994: data <= 8'h1F;
            16'd33995: data <= 8'h00;
            16'd33996: data <= 8'h1F;
            16'd33997: data <= 8'h00;
            16'd33998: data <= 8'h1F;
            16'd33999: data <= 8'h00;
            16'd34000: data <= 8'hFF;
            16'd34001: data <= 8'hFF;
            16'd34002: data <= 8'h1F;
            16'd34003: data <= 8'h00;
            16'd34004: data <= 8'h1F;
            16'd34005: data <= 8'h00;
            16'd34006: data <= 8'h1F;
            16'd34007: data <= 8'h00;
            16'd34008: data <= 8'h1F;
            16'd34009: data <= 8'h00;
            16'd34010: data <= 8'h1F;
            16'd34011: data <= 8'h00;
            16'd34012: data <= 8'h1F;
            16'd34013: data <= 8'h00;
            16'd34014: data <= 8'h1F;
            16'd34015: data <= 8'h00;
            16'd34016: data <= 8'h1F;
            16'd34017: data <= 8'h00;
            16'd34018: data <= 8'h1F;
            16'd34019: data <= 8'h00;
            16'd34020: data <= 8'h1F;
            16'd34021: data <= 8'h00;
            16'd34022: data <= 8'h1F;
            16'd34023: data <= 8'h00;
            16'd34024: data <= 8'h1F;
            16'd34025: data <= 8'h00;
            16'd34026: data <= 8'h1F;
            16'd34027: data <= 8'h00;
            16'd34028: data <= 8'h1F;
            16'd34029: data <= 8'h00;
            16'd34030: data <= 8'h1F;
            16'd34031: data <= 8'h00;
            16'd34032: data <= 8'h1F;
            16'd34033: data <= 8'h00;
            16'd34034: data <= 8'h1F;
            16'd34035: data <= 8'h00;
            16'd34036: data <= 8'h1F;
            16'd34037: data <= 8'h00;
            16'd34038: data <= 8'h1F;
            16'd34039: data <= 8'h00;
            16'd34040: data <= 8'hFF;
            16'd34041: data <= 8'hFF;
            16'd34042: data <= 8'h1F;
            16'd34043: data <= 8'h00;
            16'd34044: data <= 8'h1F;
            16'd34045: data <= 8'h00;
            16'd34046: data <= 8'h1F;
            16'd34047: data <= 8'h00;
            16'd34048: data <= 8'h1F;
            16'd34049: data <= 8'h00;
            16'd34050: data <= 8'h1F;
            16'd34051: data <= 8'h00;
            16'd34052: data <= 8'h1F;
            16'd34053: data <= 8'h00;
            16'd34054: data <= 8'h1F;
            16'd34055: data <= 8'h00;
            16'd34056: data <= 8'h1F;
            16'd34057: data <= 8'h00;
            16'd34058: data <= 8'h1F;
            16'd34059: data <= 8'h00;
            16'd34060: data <= 8'h1F;
            16'd34061: data <= 8'h00;
            16'd34062: data <= 8'h1F;
            16'd34063: data <= 8'h00;
            16'd34064: data <= 8'h1F;
            16'd34065: data <= 8'h00;
            16'd34066: data <= 8'h1F;
            16'd34067: data <= 8'h00;
            16'd34068: data <= 8'h1F;
            16'd34069: data <= 8'h00;
            16'd34070: data <= 8'h1F;
            16'd34071: data <= 8'h00;
            16'd34072: data <= 8'h1F;
            16'd34073: data <= 8'h00;
            16'd34074: data <= 8'h1F;
            16'd34075: data <= 8'h00;
            16'd34076: data <= 8'h1F;
            16'd34077: data <= 8'h00;
            16'd34078: data <= 8'h1F;
            16'd34079: data <= 8'h00;
            16'd34080: data <= 8'hFF;
            16'd34081: data <= 8'hFF;
            16'd34082: data <= 8'h1F;
            16'd34083: data <= 8'h00;
            16'd34084: data <= 8'h1F;
            16'd34085: data <= 8'h00;
            16'd34086: data <= 8'h1F;
            16'd34087: data <= 8'h00;
            16'd34088: data <= 8'h1F;
            16'd34089: data <= 8'h00;
            16'd34090: data <= 8'h1F;
            16'd34091: data <= 8'h00;
            16'd34092: data <= 8'h1F;
            16'd34093: data <= 8'h00;
            16'd34094: data <= 8'h1F;
            16'd34095: data <= 8'h00;
            16'd34096: data <= 8'h1F;
            16'd34097: data <= 8'h00;
            16'd34098: data <= 8'h1F;
            16'd34099: data <= 8'h00;
            16'd34100: data <= 8'h1F;
            16'd34101: data <= 8'h00;
            16'd34102: data <= 8'h1F;
            16'd34103: data <= 8'h00;
            16'd34104: data <= 8'h1F;
            16'd34105: data <= 8'h00;
            16'd34106: data <= 8'h1F;
            16'd34107: data <= 8'h00;
            16'd34108: data <= 8'h1F;
            16'd34109: data <= 8'h00;
            16'd34110: data <= 8'h1F;
            16'd34111: data <= 8'h00;
            16'd34112: data <= 8'h1F;
            16'd34113: data <= 8'h00;
            16'd34114: data <= 8'h1F;
            16'd34115: data <= 8'h00;
            16'd34116: data <= 8'h1F;
            16'd34117: data <= 8'h00;
            16'd34118: data <= 8'h1F;
            16'd34119: data <= 8'h00;
            16'd34120: data <= 8'hFF;
            16'd34121: data <= 8'hFF;
            16'd34122: data <= 8'h1F;
            16'd34123: data <= 8'h00;
            16'd34124: data <= 8'h1F;
            16'd34125: data <= 8'h00;
            16'd34126: data <= 8'h1F;
            16'd34127: data <= 8'h00;
            16'd34128: data <= 8'h1F;
            16'd34129: data <= 8'h00;
            16'd34130: data <= 8'h1F;
            16'd34131: data <= 8'h00;
            16'd34132: data <= 8'h1F;
            16'd34133: data <= 8'h00;
            16'd34134: data <= 8'h1F;
            16'd34135: data <= 8'h00;
            16'd34136: data <= 8'h1F;
            16'd34137: data <= 8'h00;
            16'd34138: data <= 8'h1F;
            16'd34139: data <= 8'h00;
            16'd34140: data <= 8'h1F;
            16'd34141: data <= 8'h00;
            16'd34142: data <= 8'h1F;
            16'd34143: data <= 8'h00;
            16'd34144: data <= 8'h1F;
            16'd34145: data <= 8'h00;
            16'd34146: data <= 8'h1F;
            16'd34147: data <= 8'h00;
            16'd34148: data <= 8'h1F;
            16'd34149: data <= 8'h00;
            16'd34150: data <= 8'h1F;
            16'd34151: data <= 8'h00;
            16'd34152: data <= 8'h1F;
            16'd34153: data <= 8'h00;
            16'd34154: data <= 8'h1F;
            16'd34155: data <= 8'h00;
            16'd34156: data <= 8'h1F;
            16'd34157: data <= 8'h00;
            16'd34158: data <= 8'h1F;
            16'd34159: data <= 8'h00;
            16'd34160: data <= 8'hFF;
            16'd34161: data <= 8'hFF;
            16'd34162: data <= 8'h1F;
            16'd34163: data <= 8'h00;
            16'd34164: data <= 8'h1F;
            16'd34165: data <= 8'h00;
            16'd34166: data <= 8'h1F;
            16'd34167: data <= 8'h00;
            16'd34168: data <= 8'h1F;
            16'd34169: data <= 8'h00;
            16'd34170: data <= 8'h1F;
            16'd34171: data <= 8'h00;
            16'd34172: data <= 8'h1F;
            16'd34173: data <= 8'h00;
            16'd34174: data <= 8'h1F;
            16'd34175: data <= 8'h00;
            16'd34176: data <= 8'h1F;
            16'd34177: data <= 8'h00;
            16'd34178: data <= 8'h1F;
            16'd34179: data <= 8'h00;
            16'd34180: data <= 8'h1F;
            16'd34181: data <= 8'h00;
            16'd34182: data <= 8'h1F;
            16'd34183: data <= 8'h00;
            16'd34184: data <= 8'h1F;
            16'd34185: data <= 8'h00;
            16'd34186: data <= 8'h1F;
            16'd34187: data <= 8'h00;
            16'd34188: data <= 8'h1F;
            16'd34189: data <= 8'h00;
            16'd34190: data <= 8'h1F;
            16'd34191: data <= 8'h00;
            16'd34192: data <= 8'h1F;
            16'd34193: data <= 8'h00;
            16'd34194: data <= 8'h1F;
            16'd34195: data <= 8'h00;
            16'd34196: data <= 8'h1F;
            16'd34197: data <= 8'h00;
            16'd34198: data <= 8'h1F;
            16'd34199: data <= 8'h00;
            16'd34200: data <= 8'hFF;
            16'd34201: data <= 8'hFF;
            16'd34202: data <= 8'h1F;
            16'd34203: data <= 8'h00;
            16'd34204: data <= 8'h1F;
            16'd34205: data <= 8'h00;
            16'd34206: data <= 8'h1F;
            16'd34207: data <= 8'h00;
            16'd34208: data <= 8'h1F;
            16'd34209: data <= 8'h00;
            16'd34210: data <= 8'h1F;
            16'd34211: data <= 8'h00;
            16'd34212: data <= 8'h1F;
            16'd34213: data <= 8'h00;
            16'd34214: data <= 8'h1F;
            16'd34215: data <= 8'h00;
            16'd34216: data <= 8'h1F;
            16'd34217: data <= 8'h00;
            16'd34218: data <= 8'h1F;
            16'd34219: data <= 8'h00;
            16'd34220: data <= 8'h1F;
            16'd34221: data <= 8'h00;
            16'd34222: data <= 8'h1F;
            16'd34223: data <= 8'h00;
            16'd34224: data <= 8'h1F;
            16'd34225: data <= 8'h00;
            16'd34226: data <= 8'h1F;
            16'd34227: data <= 8'h00;
            16'd34228: data <= 8'h1F;
            16'd34229: data <= 8'h00;
            16'd34230: data <= 8'h1F;
            16'd34231: data <= 8'h00;
            16'd34232: data <= 8'h1F;
            16'd34233: data <= 8'h00;
            16'd34234: data <= 8'h1F;
            16'd34235: data <= 8'h00;
            16'd34236: data <= 8'h1F;
            16'd34237: data <= 8'h00;
            16'd34238: data <= 8'h1F;
            16'd34239: data <= 8'h00;
            16'd34240: data <= 8'hFF;
            16'd34241: data <= 8'hFF;
            16'd34242: data <= 8'h1F;
            16'd34243: data <= 8'h00;
            16'd34244: data <= 8'h1F;
            16'd34245: data <= 8'h00;
            16'd34246: data <= 8'h1F;
            16'd34247: data <= 8'h00;
            16'd34248: data <= 8'h1F;
            16'd34249: data <= 8'h00;
            16'd34250: data <= 8'h1F;
            16'd34251: data <= 8'h00;
            16'd34252: data <= 8'h1F;
            16'd34253: data <= 8'h00;
            16'd34254: data <= 8'h1F;
            16'd34255: data <= 8'h00;
            16'd34256: data <= 8'h1F;
            16'd34257: data <= 8'h00;
            16'd34258: data <= 8'h1F;
            16'd34259: data <= 8'h00;
            16'd34260: data <= 8'h1F;
            16'd34261: data <= 8'h00;
            16'd34262: data <= 8'h1F;
            16'd34263: data <= 8'h00;
            16'd34264: data <= 8'h1F;
            16'd34265: data <= 8'h00;
            16'd34266: data <= 8'h1F;
            16'd34267: data <= 8'h00;
            16'd34268: data <= 8'h1F;
            16'd34269: data <= 8'h00;
            16'd34270: data <= 8'h1F;
            16'd34271: data <= 8'h00;
            16'd34272: data <= 8'h1F;
            16'd34273: data <= 8'h00;
            16'd34274: data <= 8'h1F;
            16'd34275: data <= 8'h00;
            16'd34276: data <= 8'h1F;
            16'd34277: data <= 8'h00;
            16'd34278: data <= 8'h1F;
            16'd34279: data <= 8'h00;
            16'd34280: data <= 8'hFF;
            16'd34281: data <= 8'hFF;
            16'd34282: data <= 8'h1F;
            16'd34283: data <= 8'h00;
            16'd34284: data <= 8'h1F;
            16'd34285: data <= 8'h00;
            16'd34286: data <= 8'h1F;
            16'd34287: data <= 8'h00;
            16'd34288: data <= 8'h1F;
            16'd34289: data <= 8'h00;
            16'd34290: data <= 8'h1F;
            16'd34291: data <= 8'h00;
            16'd34292: data <= 8'h1F;
            16'd34293: data <= 8'h00;
            16'd34294: data <= 8'h1F;
            16'd34295: data <= 8'h00;
            16'd34296: data <= 8'h1F;
            16'd34297: data <= 8'h00;
            16'd34298: data <= 8'h1F;
            16'd34299: data <= 8'h00;
            16'd34300: data <= 8'h1F;
            16'd34301: data <= 8'h00;
            16'd34302: data <= 8'h1F;
            16'd34303: data <= 8'h00;
            16'd34304: data <= 8'h1F;
            16'd34305: data <= 8'h00;
            16'd34306: data <= 8'h1F;
            16'd34307: data <= 8'h00;
            16'd34308: data <= 8'h1F;
            16'd34309: data <= 8'h00;
            16'd34310: data <= 8'h1F;
            16'd34311: data <= 8'h00;
            16'd34312: data <= 8'h1F;
            16'd34313: data <= 8'h00;
            16'd34314: data <= 8'h1F;
            16'd34315: data <= 8'h00;
            16'd34316: data <= 8'h1F;
            16'd34317: data <= 8'h00;
            16'd34318: data <= 8'h1F;
            16'd34319: data <= 8'h00;
            16'd34320: data <= 8'hFF;
            16'd34321: data <= 8'hFF;
            16'd34322: data <= 8'h1F;
            16'd34323: data <= 8'h00;
            16'd34324: data <= 8'h1F;
            16'd34325: data <= 8'h00;
            16'd34326: data <= 8'h1F;
            16'd34327: data <= 8'h00;
            16'd34328: data <= 8'h1F;
            16'd34329: data <= 8'h00;
            16'd34330: data <= 8'h1F;
            16'd34331: data <= 8'h00;
            16'd34332: data <= 8'h1F;
            16'd34333: data <= 8'h00;
            16'd34334: data <= 8'h1F;
            16'd34335: data <= 8'h00;
            16'd34336: data <= 8'h1F;
            16'd34337: data <= 8'h00;
            16'd34338: data <= 8'h1F;
            16'd34339: data <= 8'h00;
            16'd34340: data <= 8'h1F;
            16'd34341: data <= 8'h00;
            16'd34342: data <= 8'h1F;
            16'd34343: data <= 8'h00;
            16'd34344: data <= 8'h1F;
            16'd34345: data <= 8'h00;
            16'd34346: data <= 8'h1F;
            16'd34347: data <= 8'h00;
            16'd34348: data <= 8'h1F;
            16'd34349: data <= 8'h00;
            16'd34350: data <= 8'h1F;
            16'd34351: data <= 8'h00;
            16'd34352: data <= 8'h1F;
            16'd34353: data <= 8'h00;
            16'd34354: data <= 8'h1F;
            16'd34355: data <= 8'h00;
            16'd34356: data <= 8'h1F;
            16'd34357: data <= 8'h00;
            16'd34358: data <= 8'h1F;
            16'd34359: data <= 8'h00;
            16'd34360: data <= 8'hFF;
            16'd34361: data <= 8'hFF;
            16'd34362: data <= 8'h1F;
            16'd34363: data <= 8'h00;
            16'd34364: data <= 8'h1F;
            16'd34365: data <= 8'h00;
            16'd34366: data <= 8'h1F;
            16'd34367: data <= 8'h00;
            16'd34368: data <= 8'h1F;
            16'd34369: data <= 8'h00;
            16'd34370: data <= 8'h1F;
            16'd34371: data <= 8'h00;
            16'd34372: data <= 8'h1F;
            16'd34373: data <= 8'h00;
            16'd34374: data <= 8'h1F;
            16'd34375: data <= 8'h00;
            16'd34376: data <= 8'h1F;
            16'd34377: data <= 8'h00;
            16'd34378: data <= 8'h1F;
            16'd34379: data <= 8'h00;
            16'd34380: data <= 8'h1F;
            16'd34381: data <= 8'h00;
            16'd34382: data <= 8'h1F;
            16'd34383: data <= 8'h00;
            16'd34384: data <= 8'h1F;
            16'd34385: data <= 8'h00;
            16'd34386: data <= 8'h1F;
            16'd34387: data <= 8'h00;
            16'd34388: data <= 8'h1F;
            16'd34389: data <= 8'h00;
            16'd34390: data <= 8'h1F;
            16'd34391: data <= 8'h00;
            16'd34392: data <= 8'h1F;
            16'd34393: data <= 8'h00;
            16'd34394: data <= 8'h1F;
            16'd34395: data <= 8'h00;
            16'd34396: data <= 8'h1F;
            16'd34397: data <= 8'h00;
            16'd34398: data <= 8'h1F;
            16'd34399: data <= 8'h00;
            16'd34400: data <= 8'hFF;
            16'd34401: data <= 8'hFF;
            16'd34402: data <= 8'h1F;
            16'd34403: data <= 8'h00;
            16'd34404: data <= 8'h1F;
            16'd34405: data <= 8'h00;
            16'd34406: data <= 8'h1F;
            16'd34407: data <= 8'h00;
            16'd34408: data <= 8'h1F;
            16'd34409: data <= 8'h00;
            16'd34410: data <= 8'h1F;
            16'd34411: data <= 8'h00;
            16'd34412: data <= 8'h1F;
            16'd34413: data <= 8'h00;
            16'd34414: data <= 8'h1F;
            16'd34415: data <= 8'h00;
            16'd34416: data <= 8'h1F;
            16'd34417: data <= 8'h00;
            16'd34418: data <= 8'h1F;
            16'd34419: data <= 8'h00;
            16'd34420: data <= 8'h1F;
            16'd34421: data <= 8'h00;
            16'd34422: data <= 8'h1F;
            16'd34423: data <= 8'h00;
            16'd34424: data <= 8'h1F;
            16'd34425: data <= 8'h00;
            16'd34426: data <= 8'h1F;
            16'd34427: data <= 8'h00;
            16'd34428: data <= 8'h1F;
            16'd34429: data <= 8'h00;
            16'd34430: data <= 8'h1F;
            16'd34431: data <= 8'h00;
            16'd34432: data <= 8'h1F;
            16'd34433: data <= 8'h00;
            16'd34434: data <= 8'h1F;
            16'd34435: data <= 8'h00;
            16'd34436: data <= 8'h1F;
            16'd34437: data <= 8'h00;
            16'd34438: data <= 8'h1F;
            16'd34439: data <= 8'h00;
            16'd34440: data <= 8'hFF;
            16'd34441: data <= 8'hFF;
            16'd34442: data <= 8'h1F;
            16'd34443: data <= 8'h00;
            16'd34444: data <= 8'h1F;
            16'd34445: data <= 8'h00;
            16'd34446: data <= 8'h1F;
            16'd34447: data <= 8'h00;
            16'd34448: data <= 8'h1F;
            16'd34449: data <= 8'h00;
            16'd34450: data <= 8'h1F;
            16'd34451: data <= 8'h00;
            16'd34452: data <= 8'h1F;
            16'd34453: data <= 8'h00;
            16'd34454: data <= 8'h1F;
            16'd34455: data <= 8'h00;
            16'd34456: data <= 8'h1F;
            16'd34457: data <= 8'h00;
            16'd34458: data <= 8'h1F;
            16'd34459: data <= 8'h00;
            16'd34460: data <= 8'h1F;
            16'd34461: data <= 8'h00;
            16'd34462: data <= 8'h1F;
            16'd34463: data <= 8'h00;
            16'd34464: data <= 8'h1F;
            16'd34465: data <= 8'h00;
            16'd34466: data <= 8'h1F;
            16'd34467: data <= 8'h00;
            16'd34468: data <= 8'h1F;
            16'd34469: data <= 8'h00;
            16'd34470: data <= 8'h1F;
            16'd34471: data <= 8'h00;
            16'd34472: data <= 8'h1F;
            16'd34473: data <= 8'h00;
            16'd34474: data <= 8'h1F;
            16'd34475: data <= 8'h00;
            16'd34476: data <= 8'h1F;
            16'd34477: data <= 8'h00;
            16'd34478: data <= 8'h1F;
            16'd34479: data <= 8'h00;
            16'd34480: data <= 8'hFF;
            16'd34481: data <= 8'hFF;
            16'd34482: data <= 8'h1F;
            16'd34483: data <= 8'h00;
            16'd34484: data <= 8'h1F;
            16'd34485: data <= 8'h00;
            16'd34486: data <= 8'h1F;
            16'd34487: data <= 8'h00;
            16'd34488: data <= 8'h1F;
            16'd34489: data <= 8'h00;
            16'd34490: data <= 8'h1F;
            16'd34491: data <= 8'h00;
            16'd34492: data <= 8'h1F;
            16'd34493: data <= 8'h00;
            16'd34494: data <= 8'h1F;
            16'd34495: data <= 8'h00;
            16'd34496: data <= 8'h1F;
            16'd34497: data <= 8'h00;
            16'd34498: data <= 8'h1F;
            16'd34499: data <= 8'h00;
            16'd34500: data <= 8'h1F;
            16'd34501: data <= 8'h00;
            16'd34502: data <= 8'h1F;
            16'd34503: data <= 8'h00;
            16'd34504: data <= 8'h1F;
            16'd34505: data <= 8'h00;
            16'd34506: data <= 8'h1F;
            16'd34507: data <= 8'h00;
            16'd34508: data <= 8'h1F;
            16'd34509: data <= 8'h00;
            16'd34510: data <= 8'h1F;
            16'd34511: data <= 8'h00;
            16'd34512: data <= 8'h1F;
            16'd34513: data <= 8'h00;
            16'd34514: data <= 8'h1F;
            16'd34515: data <= 8'h00;
            16'd34516: data <= 8'h1F;
            16'd34517: data <= 8'h00;
            16'd34518: data <= 8'h1F;
            16'd34519: data <= 8'h00;
            16'd34520: data <= 8'hFF;
            16'd34521: data <= 8'hFF;
            16'd34522: data <= 8'h1F;
            16'd34523: data <= 8'h00;
            16'd34524: data <= 8'h1F;
            16'd34525: data <= 8'h00;
            16'd34526: data <= 8'h1F;
            16'd34527: data <= 8'h00;
            16'd34528: data <= 8'h1F;
            16'd34529: data <= 8'h00;
            16'd34530: data <= 8'h1F;
            16'd34531: data <= 8'h00;
            16'd34532: data <= 8'h1F;
            16'd34533: data <= 8'h00;
            16'd34534: data <= 8'h1F;
            16'd34535: data <= 8'h00;
            16'd34536: data <= 8'h1F;
            16'd34537: data <= 8'h00;
            16'd34538: data <= 8'h1F;
            16'd34539: data <= 8'h00;
            16'd34540: data <= 8'h1F;
            16'd34541: data <= 8'h00;
            16'd34542: data <= 8'h1F;
            16'd34543: data <= 8'h00;
            16'd34544: data <= 8'h1F;
            16'd34545: data <= 8'h00;
            16'd34546: data <= 8'h1F;
            16'd34547: data <= 8'h00;
            16'd34548: data <= 8'h1F;
            16'd34549: data <= 8'h00;
            16'd34550: data <= 8'h1F;
            16'd34551: data <= 8'h00;
            16'd34552: data <= 8'h1F;
            16'd34553: data <= 8'h00;
            16'd34554: data <= 8'h1F;
            16'd34555: data <= 8'h00;
            16'd34556: data <= 8'h1F;
            16'd34557: data <= 8'h00;
            16'd34558: data <= 8'h1F;
            16'd34559: data <= 8'h00;
            16'd34560: data <= 8'hFF;
            16'd34561: data <= 8'hFF;
            16'd34562: data <= 8'h1F;
            16'd34563: data <= 8'h00;
            16'd34564: data <= 8'h1F;
            16'd34565: data <= 8'h00;
            16'd34566: data <= 8'h1F;
            16'd34567: data <= 8'h00;
            16'd34568: data <= 8'h1F;
            16'd34569: data <= 8'h00;
            16'd34570: data <= 8'h1F;
            16'd34571: data <= 8'h00;
            16'd34572: data <= 8'h1F;
            16'd34573: data <= 8'h00;
            16'd34574: data <= 8'h1F;
            16'd34575: data <= 8'h00;
            16'd34576: data <= 8'h1F;
            16'd34577: data <= 8'h00;
            16'd34578: data <= 8'h1F;
            16'd34579: data <= 8'h00;
            16'd34580: data <= 8'h1F;
            16'd34581: data <= 8'h00;
            16'd34582: data <= 8'h1F;
            16'd34583: data <= 8'h00;
            16'd34584: data <= 8'h1F;
            16'd34585: data <= 8'h00;
            16'd34586: data <= 8'h1F;
            16'd34587: data <= 8'h00;
            16'd34588: data <= 8'h1F;
            16'd34589: data <= 8'h00;
            16'd34590: data <= 8'h1F;
            16'd34591: data <= 8'h00;
            16'd34592: data <= 8'h1F;
            16'd34593: data <= 8'h00;
            16'd34594: data <= 8'h1F;
            16'd34595: data <= 8'h00;
            16'd34596: data <= 8'h1F;
            16'd34597: data <= 8'h00;
            16'd34598: data <= 8'h1F;
            16'd34599: data <= 8'h00;
            16'd34600: data <= 8'hFF;
            16'd34601: data <= 8'hFF;
            16'd34602: data <= 8'h1F;
            16'd34603: data <= 8'h00;
            16'd34604: data <= 8'h1F;
            16'd34605: data <= 8'h00;
            16'd34606: data <= 8'h1F;
            16'd34607: data <= 8'h00;
            16'd34608: data <= 8'h1F;
            16'd34609: data <= 8'h00;
            16'd34610: data <= 8'h1F;
            16'd34611: data <= 8'h00;
            16'd34612: data <= 8'h1F;
            16'd34613: data <= 8'h00;
            16'd34614: data <= 8'h1F;
            16'd34615: data <= 8'h00;
            16'd34616: data <= 8'h1F;
            16'd34617: data <= 8'h00;
            16'd34618: data <= 8'h1F;
            16'd34619: data <= 8'h00;
            16'd34620: data <= 8'h1F;
            16'd34621: data <= 8'h00;
            16'd34622: data <= 8'h1F;
            16'd34623: data <= 8'h00;
            16'd34624: data <= 8'h1F;
            16'd34625: data <= 8'h00;
            16'd34626: data <= 8'h1F;
            16'd34627: data <= 8'h00;
            16'd34628: data <= 8'h1F;
            16'd34629: data <= 8'h00;
            16'd34630: data <= 8'h1F;
            16'd34631: data <= 8'h00;
            16'd34632: data <= 8'h1F;
            16'd34633: data <= 8'h00;
            16'd34634: data <= 8'h1F;
            16'd34635: data <= 8'h00;
            16'd34636: data <= 8'h1F;
            16'd34637: data <= 8'h00;
            16'd34638: data <= 8'h1F;
            16'd34639: data <= 8'h00;
            16'd34640: data <= 8'hFF;
            16'd34641: data <= 8'hFF;
            16'd34642: data <= 8'h1F;
            16'd34643: data <= 8'h00;
            16'd34644: data <= 8'h1F;
            16'd34645: data <= 8'h00;
            16'd34646: data <= 8'h1F;
            16'd34647: data <= 8'h00;
            16'd34648: data <= 8'h1F;
            16'd34649: data <= 8'h00;
            16'd34650: data <= 8'h1F;
            16'd34651: data <= 8'h00;
            16'd34652: data <= 8'h1F;
            16'd34653: data <= 8'h00;
            16'd34654: data <= 8'h1F;
            16'd34655: data <= 8'h00;
            16'd34656: data <= 8'h1F;
            16'd34657: data <= 8'h00;
            16'd34658: data <= 8'h1F;
            16'd34659: data <= 8'h00;
            16'd34660: data <= 8'h1F;
            16'd34661: data <= 8'h00;
            16'd34662: data <= 8'h1F;
            16'd34663: data <= 8'h00;
            16'd34664: data <= 8'h1F;
            16'd34665: data <= 8'h00;
            16'd34666: data <= 8'h1F;
            16'd34667: data <= 8'h00;
            16'd34668: data <= 8'h1F;
            16'd34669: data <= 8'h00;
            16'd34670: data <= 8'h1F;
            16'd34671: data <= 8'h00;
            16'd34672: data <= 8'h1F;
            16'd34673: data <= 8'h00;
            16'd34674: data <= 8'h1F;
            16'd34675: data <= 8'h00;
            16'd34676: data <= 8'h1F;
            16'd34677: data <= 8'h00;
            16'd34678: data <= 8'h1F;
            16'd34679: data <= 8'h00;
            16'd34680: data <= 8'hFF;
            16'd34681: data <= 8'hFF;
            16'd34682: data <= 8'h1F;
            16'd34683: data <= 8'h00;
            16'd34684: data <= 8'h1F;
            16'd34685: data <= 8'h00;
            16'd34686: data <= 8'h1F;
            16'd34687: data <= 8'h00;
            16'd34688: data <= 8'h1F;
            16'd34689: data <= 8'h00;
            16'd34690: data <= 8'h1F;
            16'd34691: data <= 8'h00;
            16'd34692: data <= 8'h1F;
            16'd34693: data <= 8'h00;
            16'd34694: data <= 8'h1F;
            16'd34695: data <= 8'h00;
            16'd34696: data <= 8'h1F;
            16'd34697: data <= 8'h00;
            16'd34698: data <= 8'h1F;
            16'd34699: data <= 8'h00;
            16'd34700: data <= 8'h1F;
            16'd34701: data <= 8'h00;
            16'd34702: data <= 8'h1F;
            16'd34703: data <= 8'h00;
            16'd34704: data <= 8'h1F;
            16'd34705: data <= 8'h00;
            16'd34706: data <= 8'h1F;
            16'd34707: data <= 8'h00;
            16'd34708: data <= 8'h1F;
            16'd34709: data <= 8'h00;
            16'd34710: data <= 8'h1F;
            16'd34711: data <= 8'h00;
            16'd34712: data <= 8'h1F;
            16'd34713: data <= 8'h00;
            16'd34714: data <= 8'h1F;
            16'd34715: data <= 8'h00;
            16'd34716: data <= 8'h1F;
            16'd34717: data <= 8'h00;
            16'd34718: data <= 8'h1F;
            16'd34719: data <= 8'h00;
            16'd34720: data <= 8'hFF;
            16'd34721: data <= 8'hFF;
            16'd34722: data <= 8'h1F;
            16'd34723: data <= 8'h00;
            16'd34724: data <= 8'h1F;
            16'd34725: data <= 8'h00;
            16'd34726: data <= 8'h1F;
            16'd34727: data <= 8'h00;
            16'd34728: data <= 8'h1F;
            16'd34729: data <= 8'h00;
            16'd34730: data <= 8'h1F;
            16'd34731: data <= 8'h00;
            16'd34732: data <= 8'h1F;
            16'd34733: data <= 8'h00;
            16'd34734: data <= 8'h1F;
            16'd34735: data <= 8'h00;
            16'd34736: data <= 8'h1F;
            16'd34737: data <= 8'h00;
            16'd34738: data <= 8'h1F;
            16'd34739: data <= 8'h00;
            16'd34740: data <= 8'h1F;
            16'd34741: data <= 8'h00;
            16'd34742: data <= 8'h1F;
            16'd34743: data <= 8'h00;
            16'd34744: data <= 8'h1F;
            16'd34745: data <= 8'h00;
            16'd34746: data <= 8'h1F;
            16'd34747: data <= 8'h00;
            16'd34748: data <= 8'h1F;
            16'd34749: data <= 8'h00;
            16'd34750: data <= 8'h1F;
            16'd34751: data <= 8'h00;
            16'd34752: data <= 8'h1F;
            16'd34753: data <= 8'h00;
            16'd34754: data <= 8'h1F;
            16'd34755: data <= 8'h00;
            16'd34756: data <= 8'h1F;
            16'd34757: data <= 8'h00;
            16'd34758: data <= 8'h1F;
            16'd34759: data <= 8'h00;
            16'd34760: data <= 8'hFF;
            16'd34761: data <= 8'hFF;
            16'd34762: data <= 8'h1F;
            16'd34763: data <= 8'h00;
            16'd34764: data <= 8'h1F;
            16'd34765: data <= 8'h00;
            16'd34766: data <= 8'h1F;
            16'd34767: data <= 8'h00;
            16'd34768: data <= 8'h1F;
            16'd34769: data <= 8'h00;
            16'd34770: data <= 8'h1F;
            16'd34771: data <= 8'h00;
            16'd34772: data <= 8'h1F;
            16'd34773: data <= 8'h00;
            16'd34774: data <= 8'h1F;
            16'd34775: data <= 8'h00;
            16'd34776: data <= 8'h1F;
            16'd34777: data <= 8'h00;
            16'd34778: data <= 8'h1F;
            16'd34779: data <= 8'h00;
            16'd34780: data <= 8'h1F;
            16'd34781: data <= 8'h00;
            16'd34782: data <= 8'h1F;
            16'd34783: data <= 8'h00;
            16'd34784: data <= 8'h1F;
            16'd34785: data <= 8'h00;
            16'd34786: data <= 8'h1F;
            16'd34787: data <= 8'h00;
            16'd34788: data <= 8'h1F;
            16'd34789: data <= 8'h00;
            16'd34790: data <= 8'h1F;
            16'd34791: data <= 8'h00;
            16'd34792: data <= 8'h1F;
            16'd34793: data <= 8'h00;
            16'd34794: data <= 8'h1F;
            16'd34795: data <= 8'h00;
            16'd34796: data <= 8'h1F;
            16'd34797: data <= 8'h00;
            16'd34798: data <= 8'h1F;
            16'd34799: data <= 8'h00;
            16'd34800: data <= 8'hFF;
            16'd34801: data <= 8'hFF;
            16'd34802: data <= 8'h1F;
            16'd34803: data <= 8'h00;
            16'd34804: data <= 8'h1F;
            16'd34805: data <= 8'h00;
            16'd34806: data <= 8'h1F;
            16'd34807: data <= 8'h00;
            16'd34808: data <= 8'h1F;
            16'd34809: data <= 8'h00;
            16'd34810: data <= 8'h1F;
            16'd34811: data <= 8'h00;
            16'd34812: data <= 8'h1F;
            16'd34813: data <= 8'h00;
            16'd34814: data <= 8'h1F;
            16'd34815: data <= 8'h00;
            16'd34816: data <= 8'h1F;
            16'd34817: data <= 8'h00;
            16'd34818: data <= 8'h1F;
            16'd34819: data <= 8'h00;
            16'd34820: data <= 8'h1F;
            16'd34821: data <= 8'h00;
            16'd34822: data <= 8'h1F;
            16'd34823: data <= 8'h00;
            16'd34824: data <= 8'h1F;
            16'd34825: data <= 8'h00;
            16'd34826: data <= 8'h1F;
            16'd34827: data <= 8'h00;
            16'd34828: data <= 8'h1F;
            16'd34829: data <= 8'h00;
            16'd34830: data <= 8'h1F;
            16'd34831: data <= 8'h00;
            16'd34832: data <= 8'h1F;
            16'd34833: data <= 8'h00;
            16'd34834: data <= 8'h1F;
            16'd34835: data <= 8'h00;
            16'd34836: data <= 8'h1F;
            16'd34837: data <= 8'h00;
            16'd34838: data <= 8'h1F;
            16'd34839: data <= 8'h00;
            16'd34840: data <= 8'hFF;
            16'd34841: data <= 8'hFF;
            16'd34842: data <= 8'h1F;
            16'd34843: data <= 8'h00;
            16'd34844: data <= 8'h1F;
            16'd34845: data <= 8'h00;
            16'd34846: data <= 8'h1F;
            16'd34847: data <= 8'h00;
            16'd34848: data <= 8'h1F;
            16'd34849: data <= 8'h00;
            16'd34850: data <= 8'h1F;
            16'd34851: data <= 8'h00;
            16'd34852: data <= 8'h1F;
            16'd34853: data <= 8'h00;
            16'd34854: data <= 8'h1F;
            16'd34855: data <= 8'h00;
            16'd34856: data <= 8'h1F;
            16'd34857: data <= 8'h00;
            16'd34858: data <= 8'h1F;
            16'd34859: data <= 8'h00;
            16'd34860: data <= 8'h1F;
            16'd34861: data <= 8'h00;
            16'd34862: data <= 8'h1F;
            16'd34863: data <= 8'h00;
            16'd34864: data <= 8'h1F;
            16'd34865: data <= 8'h00;
            16'd34866: data <= 8'h1F;
            16'd34867: data <= 8'h00;
            16'd34868: data <= 8'h1F;
            16'd34869: data <= 8'h00;
            16'd34870: data <= 8'h1F;
            16'd34871: data <= 8'h00;
            16'd34872: data <= 8'h1F;
            16'd34873: data <= 8'h00;
            16'd34874: data <= 8'h1F;
            16'd34875: data <= 8'h00;
            16'd34876: data <= 8'h1F;
            16'd34877: data <= 8'h00;
            16'd34878: data <= 8'h1F;
            16'd34879: data <= 8'h00;
            16'd34880: data <= 8'hFF;
            16'd34881: data <= 8'hFF;
            16'd34882: data <= 8'h1F;
            16'd34883: data <= 8'h00;
            16'd34884: data <= 8'h1F;
            16'd34885: data <= 8'h00;
            16'd34886: data <= 8'h1F;
            16'd34887: data <= 8'h00;
            16'd34888: data <= 8'h1F;
            16'd34889: data <= 8'h00;
            16'd34890: data <= 8'h1F;
            16'd34891: data <= 8'h00;
            16'd34892: data <= 8'h1F;
            16'd34893: data <= 8'h00;
            16'd34894: data <= 8'h1F;
            16'd34895: data <= 8'h00;
            16'd34896: data <= 8'h1F;
            16'd34897: data <= 8'h00;
            16'd34898: data <= 8'h1F;
            16'd34899: data <= 8'h00;
            16'd34900: data <= 8'h1F;
            16'd34901: data <= 8'h00;
            16'd34902: data <= 8'h1F;
            16'd34903: data <= 8'h00;
            16'd34904: data <= 8'h1F;
            16'd34905: data <= 8'h00;
            16'd34906: data <= 8'h1F;
            16'd34907: data <= 8'h00;
            16'd34908: data <= 8'h1F;
            16'd34909: data <= 8'h00;
            16'd34910: data <= 8'h1F;
            16'd34911: data <= 8'h00;
            16'd34912: data <= 8'h1F;
            16'd34913: data <= 8'h00;
            16'd34914: data <= 8'h1F;
            16'd34915: data <= 8'h00;
            16'd34916: data <= 8'h1F;
            16'd34917: data <= 8'h00;
            16'd34918: data <= 8'h1F;
            16'd34919: data <= 8'h00;
            16'd34920: data <= 8'hFF;
            16'd34921: data <= 8'hFF;
            16'd34922: data <= 8'h1F;
            16'd34923: data <= 8'h00;
            16'd34924: data <= 8'h1F;
            16'd34925: data <= 8'h00;
            16'd34926: data <= 8'h1F;
            16'd34927: data <= 8'h00;
            16'd34928: data <= 8'h1F;
            16'd34929: data <= 8'h00;
            16'd34930: data <= 8'h1F;
            16'd34931: data <= 8'h00;
            16'd34932: data <= 8'h1F;
            16'd34933: data <= 8'h00;
            16'd34934: data <= 8'h1F;
            16'd34935: data <= 8'h00;
            16'd34936: data <= 8'h1F;
            16'd34937: data <= 8'h00;
            16'd34938: data <= 8'h1F;
            16'd34939: data <= 8'h00;
            16'd34940: data <= 8'h1F;
            16'd34941: data <= 8'h00;
            16'd34942: data <= 8'h1F;
            16'd34943: data <= 8'h00;
            16'd34944: data <= 8'h1F;
            16'd34945: data <= 8'h00;
            16'd34946: data <= 8'h1F;
            16'd34947: data <= 8'h00;
            16'd34948: data <= 8'h1F;
            16'd34949: data <= 8'h00;
            16'd34950: data <= 8'h1F;
            16'd34951: data <= 8'h00;
            16'd34952: data <= 8'h1F;
            16'd34953: data <= 8'h00;
            16'd34954: data <= 8'h1F;
            16'd34955: data <= 8'h00;
            16'd34956: data <= 8'h1F;
            16'd34957: data <= 8'h00;
            16'd34958: data <= 8'h1F;
            16'd34959: data <= 8'h00;
            16'd34960: data <= 8'hFF;
            16'd34961: data <= 8'hFF;
            16'd34962: data <= 8'h1F;
            16'd34963: data <= 8'h00;
            16'd34964: data <= 8'h1F;
            16'd34965: data <= 8'h00;
            16'd34966: data <= 8'h1F;
            16'd34967: data <= 8'h00;
            16'd34968: data <= 8'h1F;
            16'd34969: data <= 8'h00;
            16'd34970: data <= 8'h1F;
            16'd34971: data <= 8'h00;
            16'd34972: data <= 8'h1F;
            16'd34973: data <= 8'h00;
            16'd34974: data <= 8'h1F;
            16'd34975: data <= 8'h00;
            16'd34976: data <= 8'h1F;
            16'd34977: data <= 8'h00;
            16'd34978: data <= 8'h1F;
            16'd34979: data <= 8'h00;
            16'd34980: data <= 8'h1F;
            16'd34981: data <= 8'h00;
            16'd34982: data <= 8'h1F;
            16'd34983: data <= 8'h00;
            16'd34984: data <= 8'h1F;
            16'd34985: data <= 8'h00;
            16'd34986: data <= 8'h1F;
            16'd34987: data <= 8'h00;
            16'd34988: data <= 8'h1F;
            16'd34989: data <= 8'h00;
            16'd34990: data <= 8'h1F;
            16'd34991: data <= 8'h00;
            16'd34992: data <= 8'h1F;
            16'd34993: data <= 8'h00;
            16'd34994: data <= 8'h1F;
            16'd34995: data <= 8'h00;
            16'd34996: data <= 8'h1F;
            16'd34997: data <= 8'h00;
            16'd34998: data <= 8'h1F;
            16'd34999: data <= 8'h00;
            16'd35000: data <= 8'hFF;
            16'd35001: data <= 8'hFF;
            16'd35002: data <= 8'h1F;
            16'd35003: data <= 8'h00;
            16'd35004: data <= 8'h1F;
            16'd35005: data <= 8'h00;
            16'd35006: data <= 8'h1F;
            16'd35007: data <= 8'h00;
            16'd35008: data <= 8'h1F;
            16'd35009: data <= 8'h00;
            16'd35010: data <= 8'h1F;
            16'd35011: data <= 8'h00;
            16'd35012: data <= 8'h1F;
            16'd35013: data <= 8'h00;
            16'd35014: data <= 8'h1F;
            16'd35015: data <= 8'h00;
            16'd35016: data <= 8'h1F;
            16'd35017: data <= 8'h00;
            16'd35018: data <= 8'h1F;
            16'd35019: data <= 8'h00;
            16'd35020: data <= 8'h1F;
            16'd35021: data <= 8'h00;
            16'd35022: data <= 8'h1F;
            16'd35023: data <= 8'h00;
            16'd35024: data <= 8'h1F;
            16'd35025: data <= 8'h00;
            16'd35026: data <= 8'h1F;
            16'd35027: data <= 8'h00;
            16'd35028: data <= 8'h1F;
            16'd35029: data <= 8'h00;
            16'd35030: data <= 8'h1F;
            16'd35031: data <= 8'h00;
            16'd35032: data <= 8'h1F;
            16'd35033: data <= 8'h00;
            16'd35034: data <= 8'h1F;
            16'd35035: data <= 8'h00;
            16'd35036: data <= 8'h1F;
            16'd35037: data <= 8'h00;
            16'd35038: data <= 8'h1F;
            16'd35039: data <= 8'h00;
            16'd35040: data <= 8'hFF;
            16'd35041: data <= 8'hFF;
            16'd35042: data <= 8'h1F;
            16'd35043: data <= 8'h00;
            16'd35044: data <= 8'h1F;
            16'd35045: data <= 8'h00;
            16'd35046: data <= 8'h1F;
            16'd35047: data <= 8'h00;
            16'd35048: data <= 8'h1F;
            16'd35049: data <= 8'h00;
            16'd35050: data <= 8'h1F;
            16'd35051: data <= 8'h00;
            16'd35052: data <= 8'h1F;
            16'd35053: data <= 8'h00;
            16'd35054: data <= 8'h1F;
            16'd35055: data <= 8'h00;
            16'd35056: data <= 8'h1F;
            16'd35057: data <= 8'h00;
            16'd35058: data <= 8'h1F;
            16'd35059: data <= 8'h00;
            16'd35060: data <= 8'h1F;
            16'd35061: data <= 8'h00;
            16'd35062: data <= 8'h1F;
            16'd35063: data <= 8'h00;
            16'd35064: data <= 8'h1F;
            16'd35065: data <= 8'h00;
            16'd35066: data <= 8'h1F;
            16'd35067: data <= 8'h00;
            16'd35068: data <= 8'h1F;
            16'd35069: data <= 8'h00;
            16'd35070: data <= 8'h1F;
            16'd35071: data <= 8'h00;
            16'd35072: data <= 8'h1F;
            16'd35073: data <= 8'h00;
            16'd35074: data <= 8'h1F;
            16'd35075: data <= 8'h00;
            16'd35076: data <= 8'h1F;
            16'd35077: data <= 8'h00;
            16'd35078: data <= 8'h1F;
            16'd35079: data <= 8'h00;
            16'd35080: data <= 8'hFF;
            16'd35081: data <= 8'hFF;
            16'd35082: data <= 8'h1F;
            16'd35083: data <= 8'h00;
            16'd35084: data <= 8'h1F;
            16'd35085: data <= 8'h00;
            16'd35086: data <= 8'h1F;
            16'd35087: data <= 8'h00;
            16'd35088: data <= 8'h1F;
            16'd35089: data <= 8'h00;
            16'd35090: data <= 8'h1F;
            16'd35091: data <= 8'h00;
            16'd35092: data <= 8'h1F;
            16'd35093: data <= 8'h00;
            16'd35094: data <= 8'h1F;
            16'd35095: data <= 8'h00;
            16'd35096: data <= 8'h1F;
            16'd35097: data <= 8'h00;
            16'd35098: data <= 8'h1F;
            16'd35099: data <= 8'h00;
            16'd35100: data <= 8'h1F;
            16'd35101: data <= 8'h00;
            16'd35102: data <= 8'h1F;
            16'd35103: data <= 8'h00;
            16'd35104: data <= 8'h1F;
            16'd35105: data <= 8'h00;
            16'd35106: data <= 8'h1F;
            16'd35107: data <= 8'h00;
            16'd35108: data <= 8'h1F;
            16'd35109: data <= 8'h00;
            16'd35110: data <= 8'h1F;
            16'd35111: data <= 8'h00;
            16'd35112: data <= 8'h1F;
            16'd35113: data <= 8'h00;
            16'd35114: data <= 8'h1F;
            16'd35115: data <= 8'h00;
            16'd35116: data <= 8'h1F;
            16'd35117: data <= 8'h00;
            16'd35118: data <= 8'h1F;
            16'd35119: data <= 8'h00;
            16'd35120: data <= 8'hFF;
            16'd35121: data <= 8'hFF;
            16'd35122: data <= 8'h1F;
            16'd35123: data <= 8'h00;
            16'd35124: data <= 8'h1F;
            16'd35125: data <= 8'h00;
            16'd35126: data <= 8'h1F;
            16'd35127: data <= 8'h00;
            16'd35128: data <= 8'h1F;
            16'd35129: data <= 8'h00;
            16'd35130: data <= 8'h1F;
            16'd35131: data <= 8'h00;
            16'd35132: data <= 8'h1F;
            16'd35133: data <= 8'h00;
            16'd35134: data <= 8'h1F;
            16'd35135: data <= 8'h00;
            16'd35136: data <= 8'h1F;
            16'd35137: data <= 8'h00;
            16'd35138: data <= 8'h1F;
            16'd35139: data <= 8'h00;
            16'd35140: data <= 8'h1F;
            16'd35141: data <= 8'h00;
            16'd35142: data <= 8'h1F;
            16'd35143: data <= 8'h00;
            16'd35144: data <= 8'h1F;
            16'd35145: data <= 8'h00;
            16'd35146: data <= 8'h1F;
            16'd35147: data <= 8'h00;
            16'd35148: data <= 8'h1F;
            16'd35149: data <= 8'h00;
            16'd35150: data <= 8'h1F;
            16'd35151: data <= 8'h00;
            16'd35152: data <= 8'h1F;
            16'd35153: data <= 8'h00;
            16'd35154: data <= 8'h1F;
            16'd35155: data <= 8'h00;
            16'd35156: data <= 8'h1F;
            16'd35157: data <= 8'h00;
            16'd35158: data <= 8'h1F;
            16'd35159: data <= 8'h00;
            16'd35160: data <= 8'hFF;
            16'd35161: data <= 8'hFF;
            16'd35162: data <= 8'h1F;
            16'd35163: data <= 8'h00;
            16'd35164: data <= 8'h1F;
            16'd35165: data <= 8'h00;
            16'd35166: data <= 8'h1F;
            16'd35167: data <= 8'h00;
            16'd35168: data <= 8'h1F;
            16'd35169: data <= 8'h00;
            16'd35170: data <= 8'h1F;
            16'd35171: data <= 8'h00;
            16'd35172: data <= 8'h1F;
            16'd35173: data <= 8'h00;
            16'd35174: data <= 8'h1F;
            16'd35175: data <= 8'h00;
            16'd35176: data <= 8'h1F;
            16'd35177: data <= 8'h00;
            16'd35178: data <= 8'h1F;
            16'd35179: data <= 8'h00;
            16'd35180: data <= 8'h1F;
            16'd35181: data <= 8'h00;
            16'd35182: data <= 8'h1F;
            16'd35183: data <= 8'h00;
            16'd35184: data <= 8'h1F;
            16'd35185: data <= 8'h00;
            16'd35186: data <= 8'h1F;
            16'd35187: data <= 8'h00;
            16'd35188: data <= 8'h1F;
            16'd35189: data <= 8'h00;
            16'd35190: data <= 8'h1F;
            16'd35191: data <= 8'h00;
            16'd35192: data <= 8'h1F;
            16'd35193: data <= 8'h00;
            16'd35194: data <= 8'h1F;
            16'd35195: data <= 8'h00;
            16'd35196: data <= 8'h1F;
            16'd35197: data <= 8'h00;
            16'd35198: data <= 8'h1F;
            16'd35199: data <= 8'h00;
            16'd35200: data <= 8'hFF;
            16'd35201: data <= 8'hFF;
            16'd35202: data <= 8'h1F;
            16'd35203: data <= 8'h00;
            16'd35204: data <= 8'h1F;
            16'd35205: data <= 8'h00;
            16'd35206: data <= 8'h1F;
            16'd35207: data <= 8'h00;
            16'd35208: data <= 8'h1F;
            16'd35209: data <= 8'h00;
            16'd35210: data <= 8'h1F;
            16'd35211: data <= 8'h00;
            16'd35212: data <= 8'h1F;
            16'd35213: data <= 8'h00;
            16'd35214: data <= 8'h1F;
            16'd35215: data <= 8'h00;
            16'd35216: data <= 8'h1F;
            16'd35217: data <= 8'h00;
            16'd35218: data <= 8'h1F;
            16'd35219: data <= 8'h00;
            16'd35220: data <= 8'h1F;
            16'd35221: data <= 8'h00;
            16'd35222: data <= 8'h1F;
            16'd35223: data <= 8'h00;
            16'd35224: data <= 8'h1F;
            16'd35225: data <= 8'h00;
            16'd35226: data <= 8'h1F;
            16'd35227: data <= 8'h00;
            16'd35228: data <= 8'h1F;
            16'd35229: data <= 8'h00;
            16'd35230: data <= 8'h1F;
            16'd35231: data <= 8'h00;
            16'd35232: data <= 8'h1F;
            16'd35233: data <= 8'h00;
            16'd35234: data <= 8'h1F;
            16'd35235: data <= 8'h00;
            16'd35236: data <= 8'h1F;
            16'd35237: data <= 8'h00;
            16'd35238: data <= 8'h1F;
            16'd35239: data <= 8'h00;
            16'd35240: data <= 8'hFF;
            16'd35241: data <= 8'hFF;
            16'd35242: data <= 8'h1F;
            16'd35243: data <= 8'h00;
            16'd35244: data <= 8'h1F;
            16'd35245: data <= 8'h00;
            16'd35246: data <= 8'h1F;
            16'd35247: data <= 8'h00;
            16'd35248: data <= 8'h1F;
            16'd35249: data <= 8'h00;
            16'd35250: data <= 8'h1F;
            16'd35251: data <= 8'h00;
            16'd35252: data <= 8'h1F;
            16'd35253: data <= 8'h00;
            16'd35254: data <= 8'h1F;
            16'd35255: data <= 8'h00;
            16'd35256: data <= 8'h1F;
            16'd35257: data <= 8'h00;
            16'd35258: data <= 8'h1F;
            16'd35259: data <= 8'h00;
            16'd35260: data <= 8'h1F;
            16'd35261: data <= 8'h00;
            16'd35262: data <= 8'h1F;
            16'd35263: data <= 8'h00;
            16'd35264: data <= 8'h1F;
            16'd35265: data <= 8'h00;
            16'd35266: data <= 8'h1F;
            16'd35267: data <= 8'h00;
            16'd35268: data <= 8'h1F;
            16'd35269: data <= 8'h00;
            16'd35270: data <= 8'h1F;
            16'd35271: data <= 8'h00;
            16'd35272: data <= 8'h1F;
            16'd35273: data <= 8'h00;
            16'd35274: data <= 8'h1F;
            16'd35275: data <= 8'h00;
            16'd35276: data <= 8'h1F;
            16'd35277: data <= 8'h00;
            16'd35278: data <= 8'h1F;
            16'd35279: data <= 8'h00;
            16'd35280: data <= 8'hFF;
            16'd35281: data <= 8'hFF;
            16'd35282: data <= 8'h1F;
            16'd35283: data <= 8'h00;
            16'd35284: data <= 8'h1F;
            16'd35285: data <= 8'h00;
            16'd35286: data <= 8'h1F;
            16'd35287: data <= 8'h00;
            16'd35288: data <= 8'h1F;
            16'd35289: data <= 8'h00;
            16'd35290: data <= 8'h1F;
            16'd35291: data <= 8'h00;
            16'd35292: data <= 8'h1F;
            16'd35293: data <= 8'h00;
            16'd35294: data <= 8'h1F;
            16'd35295: data <= 8'h00;
            16'd35296: data <= 8'h1F;
            16'd35297: data <= 8'h00;
            16'd35298: data <= 8'h1F;
            16'd35299: data <= 8'h00;
            16'd35300: data <= 8'h1F;
            16'd35301: data <= 8'h00;
            16'd35302: data <= 8'h1F;
            16'd35303: data <= 8'h00;
            16'd35304: data <= 8'h1F;
            16'd35305: data <= 8'h00;
            16'd35306: data <= 8'h1F;
            16'd35307: data <= 8'h00;
            16'd35308: data <= 8'h1F;
            16'd35309: data <= 8'h00;
            16'd35310: data <= 8'h1F;
            16'd35311: data <= 8'h00;
            16'd35312: data <= 8'h1F;
            16'd35313: data <= 8'h00;
            16'd35314: data <= 8'h1F;
            16'd35315: data <= 8'h00;
            16'd35316: data <= 8'h1F;
            16'd35317: data <= 8'h00;
            16'd35318: data <= 8'h1F;
            16'd35319: data <= 8'h00;
            16'd35320: data <= 8'hFF;
            16'd35321: data <= 8'hFF;
            16'd35322: data <= 8'h1F;
            16'd35323: data <= 8'h00;
            16'd35324: data <= 8'h1F;
            16'd35325: data <= 8'h00;
            16'd35326: data <= 8'h1F;
            16'd35327: data <= 8'h00;
            16'd35328: data <= 8'h1F;
            16'd35329: data <= 8'h00;
            16'd35330: data <= 8'h1F;
            16'd35331: data <= 8'h00;
            16'd35332: data <= 8'h1F;
            16'd35333: data <= 8'h00;
            16'd35334: data <= 8'h1F;
            16'd35335: data <= 8'h00;
            16'd35336: data <= 8'h1F;
            16'd35337: data <= 8'h00;
            16'd35338: data <= 8'h1F;
            16'd35339: data <= 8'h00;
            16'd35340: data <= 8'h1F;
            16'd35341: data <= 8'h00;
            16'd35342: data <= 8'h1F;
            16'd35343: data <= 8'h00;
            16'd35344: data <= 8'h1F;
            16'd35345: data <= 8'h00;
            16'd35346: data <= 8'h1F;
            16'd35347: data <= 8'h00;
            16'd35348: data <= 8'h1F;
            16'd35349: data <= 8'h00;
            16'd35350: data <= 8'h1F;
            16'd35351: data <= 8'h00;
            16'd35352: data <= 8'h1F;
            16'd35353: data <= 8'h00;
            16'd35354: data <= 8'h1F;
            16'd35355: data <= 8'h00;
            16'd35356: data <= 8'h1F;
            16'd35357: data <= 8'h00;
            16'd35358: data <= 8'h1F;
            16'd35359: data <= 8'h00;
            16'd35360: data <= 8'hFF;
            16'd35361: data <= 8'hFF;
            16'd35362: data <= 8'h1F;
            16'd35363: data <= 8'h00;
            16'd35364: data <= 8'h1F;
            16'd35365: data <= 8'h00;
            16'd35366: data <= 8'h1F;
            16'd35367: data <= 8'h00;
            16'd35368: data <= 8'h1F;
            16'd35369: data <= 8'h00;
            16'd35370: data <= 8'h1F;
            16'd35371: data <= 8'h00;
            16'd35372: data <= 8'h1F;
            16'd35373: data <= 8'h00;
            16'd35374: data <= 8'h1F;
            16'd35375: data <= 8'h00;
            16'd35376: data <= 8'h1F;
            16'd35377: data <= 8'h00;
            16'd35378: data <= 8'h1F;
            16'd35379: data <= 8'h00;
            16'd35380: data <= 8'h1F;
            16'd35381: data <= 8'h00;
            16'd35382: data <= 8'h1F;
            16'd35383: data <= 8'h00;
            16'd35384: data <= 8'h1F;
            16'd35385: data <= 8'h00;
            16'd35386: data <= 8'h1F;
            16'd35387: data <= 8'h00;
            16'd35388: data <= 8'h1F;
            16'd35389: data <= 8'h00;
            16'd35390: data <= 8'h1F;
            16'd35391: data <= 8'h00;
            16'd35392: data <= 8'h1F;
            16'd35393: data <= 8'h00;
            16'd35394: data <= 8'h1F;
            16'd35395: data <= 8'h00;
            16'd35396: data <= 8'h1F;
            16'd35397: data <= 8'h00;
            16'd35398: data <= 8'h1F;
            16'd35399: data <= 8'h00;
            16'd35400: data <= 8'hFF;
            16'd35401: data <= 8'hFF;
            16'd35402: data <= 8'h1F;
            16'd35403: data <= 8'h00;
            16'd35404: data <= 8'h1F;
            16'd35405: data <= 8'h00;
            16'd35406: data <= 8'h1F;
            16'd35407: data <= 8'h00;
            16'd35408: data <= 8'h1F;
            16'd35409: data <= 8'h00;
            16'd35410: data <= 8'h1F;
            16'd35411: data <= 8'h00;
            16'd35412: data <= 8'h1F;
            16'd35413: data <= 8'h00;
            16'd35414: data <= 8'h1F;
            16'd35415: data <= 8'h00;
            16'd35416: data <= 8'h1F;
            16'd35417: data <= 8'h00;
            16'd35418: data <= 8'h1F;
            16'd35419: data <= 8'h00;
            16'd35420: data <= 8'h1F;
            16'd35421: data <= 8'h00;
            16'd35422: data <= 8'h1F;
            16'd35423: data <= 8'h00;
            16'd35424: data <= 8'h1F;
            16'd35425: data <= 8'h00;
            16'd35426: data <= 8'h1F;
            16'd35427: data <= 8'h00;
            16'd35428: data <= 8'h1F;
            16'd35429: data <= 8'h00;
            16'd35430: data <= 8'h1F;
            16'd35431: data <= 8'h00;
            16'd35432: data <= 8'h1F;
            16'd35433: data <= 8'h00;
            16'd35434: data <= 8'h1F;
            16'd35435: data <= 8'h00;
            16'd35436: data <= 8'h1F;
            16'd35437: data <= 8'h00;
            16'd35438: data <= 8'h1F;
            16'd35439: data <= 8'h00;
            16'd35440: data <= 8'hFF;
            16'd35441: data <= 8'hFF;
            16'd35442: data <= 8'h1F;
            16'd35443: data <= 8'h00;
            16'd35444: data <= 8'h1F;
            16'd35445: data <= 8'h00;
            16'd35446: data <= 8'h1F;
            16'd35447: data <= 8'h00;
            16'd35448: data <= 8'h1F;
            16'd35449: data <= 8'h00;
            16'd35450: data <= 8'h1F;
            16'd35451: data <= 8'h00;
            16'd35452: data <= 8'h1F;
            16'd35453: data <= 8'h00;
            16'd35454: data <= 8'h1F;
            16'd35455: data <= 8'h00;
            16'd35456: data <= 8'h1F;
            16'd35457: data <= 8'h00;
            16'd35458: data <= 8'h1F;
            16'd35459: data <= 8'h00;
            16'd35460: data <= 8'h1F;
            16'd35461: data <= 8'h00;
            16'd35462: data <= 8'h1F;
            16'd35463: data <= 8'h00;
            16'd35464: data <= 8'h1F;
            16'd35465: data <= 8'h00;
            16'd35466: data <= 8'h1F;
            16'd35467: data <= 8'h00;
            16'd35468: data <= 8'h1F;
            16'd35469: data <= 8'h00;
            16'd35470: data <= 8'h1F;
            16'd35471: data <= 8'h00;
            16'd35472: data <= 8'h1F;
            16'd35473: data <= 8'h00;
            16'd35474: data <= 8'h1F;
            16'd35475: data <= 8'h00;
            16'd35476: data <= 8'h1F;
            16'd35477: data <= 8'h00;
            16'd35478: data <= 8'h1F;
            16'd35479: data <= 8'h00;
            16'd35480: data <= 8'hFF;
            16'd35481: data <= 8'hFF;
            16'd35482: data <= 8'h1F;
            16'd35483: data <= 8'h00;
            16'd35484: data <= 8'h1F;
            16'd35485: data <= 8'h00;
            16'd35486: data <= 8'h1F;
            16'd35487: data <= 8'h00;
            16'd35488: data <= 8'h1F;
            16'd35489: data <= 8'h00;
            16'd35490: data <= 8'h1F;
            16'd35491: data <= 8'h00;
            16'd35492: data <= 8'h1F;
            16'd35493: data <= 8'h00;
            16'd35494: data <= 8'h1F;
            16'd35495: data <= 8'h00;
            16'd35496: data <= 8'h1F;
            16'd35497: data <= 8'h00;
            16'd35498: data <= 8'h1F;
            16'd35499: data <= 8'h00;
            16'd35500: data <= 8'h1F;
            16'd35501: data <= 8'h00;
            16'd35502: data <= 8'h1F;
            16'd35503: data <= 8'h00;
            16'd35504: data <= 8'h1F;
            16'd35505: data <= 8'h00;
            16'd35506: data <= 8'h1F;
            16'd35507: data <= 8'h00;
            16'd35508: data <= 8'h1F;
            16'd35509: data <= 8'h00;
            16'd35510: data <= 8'h1F;
            16'd35511: data <= 8'h00;
            16'd35512: data <= 8'h1F;
            16'd35513: data <= 8'h00;
            16'd35514: data <= 8'h1F;
            16'd35515: data <= 8'h00;
            16'd35516: data <= 8'h1F;
            16'd35517: data <= 8'h00;
            16'd35518: data <= 8'h1F;
            16'd35519: data <= 8'h00;
            16'd35520: data <= 8'hFF;
            16'd35521: data <= 8'hFF;
            16'd35522: data <= 8'h1F;
            16'd35523: data <= 8'h00;
            16'd35524: data <= 8'h1F;
            16'd35525: data <= 8'h00;
            16'd35526: data <= 8'h1F;
            16'd35527: data <= 8'h00;
            16'd35528: data <= 8'h1F;
            16'd35529: data <= 8'h00;
            16'd35530: data <= 8'h1F;
            16'd35531: data <= 8'h00;
            16'd35532: data <= 8'h1F;
            16'd35533: data <= 8'h00;
            16'd35534: data <= 8'h1F;
            16'd35535: data <= 8'h00;
            16'd35536: data <= 8'h1F;
            16'd35537: data <= 8'h00;
            16'd35538: data <= 8'h1F;
            16'd35539: data <= 8'h00;
            16'd35540: data <= 8'h1F;
            16'd35541: data <= 8'h00;
            16'd35542: data <= 8'h1F;
            16'd35543: data <= 8'h00;
            16'd35544: data <= 8'h1F;
            16'd35545: data <= 8'h00;
            16'd35546: data <= 8'h1F;
            16'd35547: data <= 8'h00;
            16'd35548: data <= 8'h1F;
            16'd35549: data <= 8'h00;
            16'd35550: data <= 8'h1F;
            16'd35551: data <= 8'h00;
            16'd35552: data <= 8'h1F;
            16'd35553: data <= 8'h00;
            16'd35554: data <= 8'h1F;
            16'd35555: data <= 8'h00;
            16'd35556: data <= 8'h1F;
            16'd35557: data <= 8'h00;
            16'd35558: data <= 8'h1F;
            16'd35559: data <= 8'h00;
            16'd35560: data <= 8'hFF;
            16'd35561: data <= 8'hFF;
            16'd35562: data <= 8'h1F;
            16'd35563: data <= 8'h00;
            16'd35564: data <= 8'h1F;
            16'd35565: data <= 8'h00;
            16'd35566: data <= 8'h1F;
            16'd35567: data <= 8'h00;
            16'd35568: data <= 8'h1F;
            16'd35569: data <= 8'h00;
            16'd35570: data <= 8'h1F;
            16'd35571: data <= 8'h00;
            16'd35572: data <= 8'h1F;
            16'd35573: data <= 8'h00;
            16'd35574: data <= 8'h1F;
            16'd35575: data <= 8'h00;
            16'd35576: data <= 8'h1F;
            16'd35577: data <= 8'h00;
            16'd35578: data <= 8'h1F;
            16'd35579: data <= 8'h00;
            16'd35580: data <= 8'h1F;
            16'd35581: data <= 8'h00;
            16'd35582: data <= 8'h1F;
            16'd35583: data <= 8'h00;
            16'd35584: data <= 8'h1F;
            16'd35585: data <= 8'h00;
            16'd35586: data <= 8'h1F;
            16'd35587: data <= 8'h00;
            16'd35588: data <= 8'h1F;
            16'd35589: data <= 8'h00;
            16'd35590: data <= 8'h1F;
            16'd35591: data <= 8'h00;
            16'd35592: data <= 8'h1F;
            16'd35593: data <= 8'h00;
            16'd35594: data <= 8'h1F;
            16'd35595: data <= 8'h00;
            16'd35596: data <= 8'h1F;
            16'd35597: data <= 8'h00;
            16'd35598: data <= 8'h1F;
            16'd35599: data <= 8'h00;
            16'd35600: data <= 8'hFF;
            16'd35601: data <= 8'hFF;
            16'd35602: data <= 8'h1F;
            16'd35603: data <= 8'h00;
            16'd35604: data <= 8'h1F;
            16'd35605: data <= 8'h00;
            16'd35606: data <= 8'h1F;
            16'd35607: data <= 8'h00;
            16'd35608: data <= 8'h1F;
            16'd35609: data <= 8'h00;
            16'd35610: data <= 8'h1F;
            16'd35611: data <= 8'h00;
            16'd35612: data <= 8'h1F;
            16'd35613: data <= 8'h00;
            16'd35614: data <= 8'h1F;
            16'd35615: data <= 8'h00;
            16'd35616: data <= 8'h1F;
            16'd35617: data <= 8'h00;
            16'd35618: data <= 8'h1F;
            16'd35619: data <= 8'h00;
            16'd35620: data <= 8'h1F;
            16'd35621: data <= 8'h00;
            16'd35622: data <= 8'h1F;
            16'd35623: data <= 8'h00;
            16'd35624: data <= 8'h1F;
            16'd35625: data <= 8'h00;
            16'd35626: data <= 8'h1F;
            16'd35627: data <= 8'h00;
            16'd35628: data <= 8'h1F;
            16'd35629: data <= 8'h00;
            16'd35630: data <= 8'h1F;
            16'd35631: data <= 8'h00;
            16'd35632: data <= 8'h1F;
            16'd35633: data <= 8'h00;
            16'd35634: data <= 8'h1F;
            16'd35635: data <= 8'h00;
            16'd35636: data <= 8'h1F;
            16'd35637: data <= 8'h00;
            16'd35638: data <= 8'h1F;
            16'd35639: data <= 8'h00;
            16'd35640: data <= 8'hFF;
            16'd35641: data <= 8'hFF;
            16'd35642: data <= 8'h1F;
            16'd35643: data <= 8'h00;
            16'd35644: data <= 8'h1F;
            16'd35645: data <= 8'h00;
            16'd35646: data <= 8'h1F;
            16'd35647: data <= 8'h00;
            16'd35648: data <= 8'h1F;
            16'd35649: data <= 8'h00;
            16'd35650: data <= 8'h1F;
            16'd35651: data <= 8'h00;
            16'd35652: data <= 8'h1F;
            16'd35653: data <= 8'h00;
            16'd35654: data <= 8'h1F;
            16'd35655: data <= 8'h00;
            16'd35656: data <= 8'h1F;
            16'd35657: data <= 8'h00;
            16'd35658: data <= 8'h1F;
            16'd35659: data <= 8'h00;
            16'd35660: data <= 8'h1F;
            16'd35661: data <= 8'h00;
            16'd35662: data <= 8'h1F;
            16'd35663: data <= 8'h00;
            16'd35664: data <= 8'h1F;
            16'd35665: data <= 8'h00;
            16'd35666: data <= 8'h1F;
            16'd35667: data <= 8'h00;
            16'd35668: data <= 8'h1F;
            16'd35669: data <= 8'h00;
            16'd35670: data <= 8'h1F;
            16'd35671: data <= 8'h00;
            16'd35672: data <= 8'h1F;
            16'd35673: data <= 8'h00;
            16'd35674: data <= 8'h1F;
            16'd35675: data <= 8'h00;
            16'd35676: data <= 8'h1F;
            16'd35677: data <= 8'h00;
            16'd35678: data <= 8'h1F;
            16'd35679: data <= 8'h00;
            16'd35680: data <= 8'hFF;
            16'd35681: data <= 8'hFF;
            16'd35682: data <= 8'h1F;
            16'd35683: data <= 8'h00;
            16'd35684: data <= 8'h1F;
            16'd35685: data <= 8'h00;
            16'd35686: data <= 8'h1F;
            16'd35687: data <= 8'h00;
            16'd35688: data <= 8'h1F;
            16'd35689: data <= 8'h00;
            16'd35690: data <= 8'h1F;
            16'd35691: data <= 8'h00;
            16'd35692: data <= 8'h1F;
            16'd35693: data <= 8'h00;
            16'd35694: data <= 8'h1F;
            16'd35695: data <= 8'h00;
            16'd35696: data <= 8'h1F;
            16'd35697: data <= 8'h00;
            16'd35698: data <= 8'h1F;
            16'd35699: data <= 8'h00;
            16'd35700: data <= 8'h1F;
            16'd35701: data <= 8'h00;
            16'd35702: data <= 8'h1F;
            16'd35703: data <= 8'h00;
            16'd35704: data <= 8'h1F;
            16'd35705: data <= 8'h00;
            16'd35706: data <= 8'h1F;
            16'd35707: data <= 8'h00;
            16'd35708: data <= 8'h1F;
            16'd35709: data <= 8'h00;
            16'd35710: data <= 8'h1F;
            16'd35711: data <= 8'h00;
            16'd35712: data <= 8'h1F;
            16'd35713: data <= 8'h00;
            16'd35714: data <= 8'h1F;
            16'd35715: data <= 8'h00;
            16'd35716: data <= 8'h1F;
            16'd35717: data <= 8'h00;
            16'd35718: data <= 8'h1F;
            16'd35719: data <= 8'h00;
            16'd35720: data <= 8'hFF;
            16'd35721: data <= 8'hFF;
            16'd35722: data <= 8'h1F;
            16'd35723: data <= 8'h00;
            16'd35724: data <= 8'h1F;
            16'd35725: data <= 8'h00;
            16'd35726: data <= 8'h1F;
            16'd35727: data <= 8'h00;
            16'd35728: data <= 8'h1F;
            16'd35729: data <= 8'h00;
            16'd35730: data <= 8'h1F;
            16'd35731: data <= 8'h00;
            16'd35732: data <= 8'h1F;
            16'd35733: data <= 8'h00;
            16'd35734: data <= 8'h1F;
            16'd35735: data <= 8'h00;
            16'd35736: data <= 8'h1F;
            16'd35737: data <= 8'h00;
            16'd35738: data <= 8'h1F;
            16'd35739: data <= 8'h00;
            16'd35740: data <= 8'h1F;
            16'd35741: data <= 8'h00;
            16'd35742: data <= 8'h1F;
            16'd35743: data <= 8'h00;
            16'd35744: data <= 8'h1F;
            16'd35745: data <= 8'h00;
            16'd35746: data <= 8'h1F;
            16'd35747: data <= 8'h00;
            16'd35748: data <= 8'h1F;
            16'd35749: data <= 8'h00;
            16'd35750: data <= 8'h1F;
            16'd35751: data <= 8'h00;
            16'd35752: data <= 8'h1F;
            16'd35753: data <= 8'h00;
            16'd35754: data <= 8'h1F;
            16'd35755: data <= 8'h00;
            16'd35756: data <= 8'h1F;
            16'd35757: data <= 8'h00;
            16'd35758: data <= 8'h1F;
            16'd35759: data <= 8'h00;
            16'd35760: data <= 8'hFF;
            16'd35761: data <= 8'hFF;
            16'd35762: data <= 8'h1F;
            16'd35763: data <= 8'h00;
            16'd35764: data <= 8'h1F;
            16'd35765: data <= 8'h00;
            16'd35766: data <= 8'h1F;
            16'd35767: data <= 8'h00;
            16'd35768: data <= 8'h1F;
            16'd35769: data <= 8'h00;
            16'd35770: data <= 8'h1F;
            16'd35771: data <= 8'h00;
            16'd35772: data <= 8'h1F;
            16'd35773: data <= 8'h00;
            16'd35774: data <= 8'h1F;
            16'd35775: data <= 8'h00;
            16'd35776: data <= 8'h1F;
            16'd35777: data <= 8'h00;
            16'd35778: data <= 8'h1F;
            16'd35779: data <= 8'h00;
            16'd35780: data <= 8'h1F;
            16'd35781: data <= 8'h00;
            16'd35782: data <= 8'h1F;
            16'd35783: data <= 8'h00;
            16'd35784: data <= 8'h1F;
            16'd35785: data <= 8'h00;
            16'd35786: data <= 8'h1F;
            16'd35787: data <= 8'h00;
            16'd35788: data <= 8'h1F;
            16'd35789: data <= 8'h00;
            16'd35790: data <= 8'h1F;
            16'd35791: data <= 8'h00;
            16'd35792: data <= 8'h1F;
            16'd35793: data <= 8'h00;
            16'd35794: data <= 8'h1F;
            16'd35795: data <= 8'h00;
            16'd35796: data <= 8'h1F;
            16'd35797: data <= 8'h00;
            16'd35798: data <= 8'h1F;
            16'd35799: data <= 8'h00;
            16'd35800: data <= 8'hFF;
            16'd35801: data <= 8'hFF;
            16'd35802: data <= 8'h1F;
            16'd35803: data <= 8'h00;
            16'd35804: data <= 8'h1F;
            16'd35805: data <= 8'h00;
            16'd35806: data <= 8'h1F;
            16'd35807: data <= 8'h00;
            16'd35808: data <= 8'h1F;
            16'd35809: data <= 8'h00;
            16'd35810: data <= 8'h1F;
            16'd35811: data <= 8'h00;
            16'd35812: data <= 8'h1F;
            16'd35813: data <= 8'h00;
            16'd35814: data <= 8'h1F;
            16'd35815: data <= 8'h00;
            16'd35816: data <= 8'h1F;
            16'd35817: data <= 8'h00;
            16'd35818: data <= 8'h1F;
            16'd35819: data <= 8'h00;
            16'd35820: data <= 8'h1F;
            16'd35821: data <= 8'h00;
            16'd35822: data <= 8'h1F;
            16'd35823: data <= 8'h00;
            16'd35824: data <= 8'h1F;
            16'd35825: data <= 8'h00;
            16'd35826: data <= 8'h1F;
            16'd35827: data <= 8'h00;
            16'd35828: data <= 8'h1F;
            16'd35829: data <= 8'h00;
            16'd35830: data <= 8'h1F;
            16'd35831: data <= 8'h00;
            16'd35832: data <= 8'h1F;
            16'd35833: data <= 8'h00;
            16'd35834: data <= 8'h1F;
            16'd35835: data <= 8'h00;
            16'd35836: data <= 8'h1F;
            16'd35837: data <= 8'h00;
            16'd35838: data <= 8'h1F;
            16'd35839: data <= 8'h00;
            16'd35840: data <= 8'hFF;
            16'd35841: data <= 8'hFF;
            16'd35842: data <= 8'h1F;
            16'd35843: data <= 8'h00;
            16'd35844: data <= 8'h1F;
            16'd35845: data <= 8'h00;
            16'd35846: data <= 8'h1F;
            16'd35847: data <= 8'h00;
            16'd35848: data <= 8'h1F;
            16'd35849: data <= 8'h00;
            16'd35850: data <= 8'h1F;
            16'd35851: data <= 8'h00;
            16'd35852: data <= 8'h1F;
            16'd35853: data <= 8'h00;
            16'd35854: data <= 8'h1F;
            16'd35855: data <= 8'h00;
            16'd35856: data <= 8'h1F;
            16'd35857: data <= 8'h00;
            16'd35858: data <= 8'h1F;
            16'd35859: data <= 8'h00;
            16'd35860: data <= 8'h1F;
            16'd35861: data <= 8'h00;
            16'd35862: data <= 8'h1F;
            16'd35863: data <= 8'h00;
            16'd35864: data <= 8'h1F;
            16'd35865: data <= 8'h00;
            16'd35866: data <= 8'h1F;
            16'd35867: data <= 8'h00;
            16'd35868: data <= 8'h1F;
            16'd35869: data <= 8'h00;
            16'd35870: data <= 8'h1F;
            16'd35871: data <= 8'h00;
            16'd35872: data <= 8'h1F;
            16'd35873: data <= 8'h00;
            16'd35874: data <= 8'h1F;
            16'd35875: data <= 8'h00;
            16'd35876: data <= 8'h1F;
            16'd35877: data <= 8'h00;
            16'd35878: data <= 8'h1F;
            16'd35879: data <= 8'h00;
            16'd35880: data <= 8'hFF;
            16'd35881: data <= 8'hFF;
            16'd35882: data <= 8'h1F;
            16'd35883: data <= 8'h00;
            16'd35884: data <= 8'h1F;
            16'd35885: data <= 8'h00;
            16'd35886: data <= 8'h1F;
            16'd35887: data <= 8'h00;
            16'd35888: data <= 8'h1F;
            16'd35889: data <= 8'h00;
            16'd35890: data <= 8'h1F;
            16'd35891: data <= 8'h00;
            16'd35892: data <= 8'h1F;
            16'd35893: data <= 8'h00;
            16'd35894: data <= 8'h1F;
            16'd35895: data <= 8'h00;
            16'd35896: data <= 8'h1F;
            16'd35897: data <= 8'h00;
            16'd35898: data <= 8'h1F;
            16'd35899: data <= 8'h00;
            16'd35900: data <= 8'h1F;
            16'd35901: data <= 8'h00;
            16'd35902: data <= 8'h1F;
            16'd35903: data <= 8'h00;
            16'd35904: data <= 8'h1F;
            16'd35905: data <= 8'h00;
            16'd35906: data <= 8'h1F;
            16'd35907: data <= 8'h00;
            16'd35908: data <= 8'h1F;
            16'd35909: data <= 8'h00;
            16'd35910: data <= 8'h1F;
            16'd35911: data <= 8'h00;
            16'd35912: data <= 8'h1F;
            16'd35913: data <= 8'h00;
            16'd35914: data <= 8'h1F;
            16'd35915: data <= 8'h00;
            16'd35916: data <= 8'h1F;
            16'd35917: data <= 8'h00;
            16'd35918: data <= 8'h1F;
            16'd35919: data <= 8'h00;
            16'd35920: data <= 8'hFF;
            16'd35921: data <= 8'hFF;
            16'd35922: data <= 8'h1F;
            16'd35923: data <= 8'h00;
            16'd35924: data <= 8'h1F;
            16'd35925: data <= 8'h00;
            16'd35926: data <= 8'h1F;
            16'd35927: data <= 8'h00;
            16'd35928: data <= 8'h1F;
            16'd35929: data <= 8'h00;
            16'd35930: data <= 8'h1F;
            16'd35931: data <= 8'h00;
            16'd35932: data <= 8'h1F;
            16'd35933: data <= 8'h00;
            16'd35934: data <= 8'h1F;
            16'd35935: data <= 8'h00;
            16'd35936: data <= 8'h1F;
            16'd35937: data <= 8'h00;
            16'd35938: data <= 8'h1F;
            16'd35939: data <= 8'h00;
            16'd35940: data <= 8'h1F;
            16'd35941: data <= 8'h00;
            16'd35942: data <= 8'h1F;
            16'd35943: data <= 8'h00;
            16'd35944: data <= 8'h1F;
            16'd35945: data <= 8'h00;
            16'd35946: data <= 8'h1F;
            16'd35947: data <= 8'h00;
            16'd35948: data <= 8'h1F;
            16'd35949: data <= 8'h00;
            16'd35950: data <= 8'h1F;
            16'd35951: data <= 8'h00;
            16'd35952: data <= 8'h1F;
            16'd35953: data <= 8'h00;
            16'd35954: data <= 8'h1F;
            16'd35955: data <= 8'h00;
            16'd35956: data <= 8'h1F;
            16'd35957: data <= 8'h00;
            16'd35958: data <= 8'h1F;
            16'd35959: data <= 8'h00;
            16'd35960: data <= 8'hFF;
            16'd35961: data <= 8'hFF;
            16'd35962: data <= 8'h1F;
            16'd35963: data <= 8'h00;
            16'd35964: data <= 8'h1F;
            16'd35965: data <= 8'h00;
            16'd35966: data <= 8'h1F;
            16'd35967: data <= 8'h00;
            16'd35968: data <= 8'h1F;
            16'd35969: data <= 8'h00;
            16'd35970: data <= 8'h1F;
            16'd35971: data <= 8'h00;
            16'd35972: data <= 8'h1F;
            16'd35973: data <= 8'h00;
            16'd35974: data <= 8'h1F;
            16'd35975: data <= 8'h00;
            16'd35976: data <= 8'h1F;
            16'd35977: data <= 8'h00;
            16'd35978: data <= 8'h1F;
            16'd35979: data <= 8'h00;
            16'd35980: data <= 8'h1F;
            16'd35981: data <= 8'h00;
            16'd35982: data <= 8'h1F;
            16'd35983: data <= 8'h00;
            16'd35984: data <= 8'h1F;
            16'd35985: data <= 8'h00;
            16'd35986: data <= 8'h1F;
            16'd35987: data <= 8'h00;
            16'd35988: data <= 8'h1F;
            16'd35989: data <= 8'h00;
            16'd35990: data <= 8'h1F;
            16'd35991: data <= 8'h00;
            16'd35992: data <= 8'h1F;
            16'd35993: data <= 8'h00;
            16'd35994: data <= 8'h1F;
            16'd35995: data <= 8'h00;
            16'd35996: data <= 8'h1F;
            16'd35997: data <= 8'h00;
            16'd35998: data <= 8'h1F;
            16'd35999: data <= 8'h00;
            16'd36000: data <= 8'hFF;
            16'd36001: data <= 8'hFF;
            16'd36002: data <= 8'h1F;
            16'd36003: data <= 8'h00;
            16'd36004: data <= 8'h1F;
            16'd36005: data <= 8'h00;
            16'd36006: data <= 8'h1F;
            16'd36007: data <= 8'h00;
            16'd36008: data <= 8'h1F;
            16'd36009: data <= 8'h00;
            16'd36010: data <= 8'h1F;
            16'd36011: data <= 8'h00;
            16'd36012: data <= 8'h1F;
            16'd36013: data <= 8'h00;
            16'd36014: data <= 8'h1F;
            16'd36015: data <= 8'h00;
            16'd36016: data <= 8'h1F;
            16'd36017: data <= 8'h00;
            16'd36018: data <= 8'h1F;
            16'd36019: data <= 8'h00;
            16'd36020: data <= 8'h1F;
            16'd36021: data <= 8'h00;
            16'd36022: data <= 8'h1F;
            16'd36023: data <= 8'h00;
            16'd36024: data <= 8'h1F;
            16'd36025: data <= 8'h00;
            16'd36026: data <= 8'h1F;
            16'd36027: data <= 8'h00;
            16'd36028: data <= 8'h1F;
            16'd36029: data <= 8'h00;
            16'd36030: data <= 8'h1F;
            16'd36031: data <= 8'h00;
            16'd36032: data <= 8'h1F;
            16'd36033: data <= 8'h00;
            16'd36034: data <= 8'h1F;
            16'd36035: data <= 8'h00;
            16'd36036: data <= 8'h1F;
            16'd36037: data <= 8'h00;
            16'd36038: data <= 8'h1F;
            16'd36039: data <= 8'h00;
            16'd36040: data <= 8'hFF;
            16'd36041: data <= 8'hFF;
            16'd36042: data <= 8'h1F;
            16'd36043: data <= 8'h00;
            16'd36044: data <= 8'h1F;
            16'd36045: data <= 8'h00;
            16'd36046: data <= 8'h1F;
            16'd36047: data <= 8'h00;
            16'd36048: data <= 8'h1F;
            16'd36049: data <= 8'h00;
            16'd36050: data <= 8'h1F;
            16'd36051: data <= 8'h00;
            16'd36052: data <= 8'h1F;
            16'd36053: data <= 8'h00;
            16'd36054: data <= 8'h1F;
            16'd36055: data <= 8'h00;
            16'd36056: data <= 8'h1F;
            16'd36057: data <= 8'h00;
            16'd36058: data <= 8'h1F;
            16'd36059: data <= 8'h00;
            16'd36060: data <= 8'h1F;
            16'd36061: data <= 8'h00;
            16'd36062: data <= 8'h1F;
            16'd36063: data <= 8'h00;
            16'd36064: data <= 8'h1F;
            16'd36065: data <= 8'h00;
            16'd36066: data <= 8'h1F;
            16'd36067: data <= 8'h00;
            16'd36068: data <= 8'h1F;
            16'd36069: data <= 8'h00;
            16'd36070: data <= 8'h1F;
            16'd36071: data <= 8'h00;
            16'd36072: data <= 8'h1F;
            16'd36073: data <= 8'h00;
            16'd36074: data <= 8'h1F;
            16'd36075: data <= 8'h00;
            16'd36076: data <= 8'h1F;
            16'd36077: data <= 8'h00;
            16'd36078: data <= 8'h1F;
            16'd36079: data <= 8'h00;
            16'd36080: data <= 8'hFF;
            16'd36081: data <= 8'hFF;
            16'd36082: data <= 8'h1F;
            16'd36083: data <= 8'h00;
            16'd36084: data <= 8'h1F;
            16'd36085: data <= 8'h00;
            16'd36086: data <= 8'h1F;
            16'd36087: data <= 8'h00;
            16'd36088: data <= 8'h1F;
            16'd36089: data <= 8'h00;
            16'd36090: data <= 8'h1F;
            16'd36091: data <= 8'h00;
            16'd36092: data <= 8'h1F;
            16'd36093: data <= 8'h00;
            16'd36094: data <= 8'h1F;
            16'd36095: data <= 8'h00;
            16'd36096: data <= 8'h1F;
            16'd36097: data <= 8'h00;
            16'd36098: data <= 8'h1F;
            16'd36099: data <= 8'h00;
            16'd36100: data <= 8'h1F;
            16'd36101: data <= 8'h00;
            16'd36102: data <= 8'h1F;
            16'd36103: data <= 8'h00;
            16'd36104: data <= 8'h1F;
            16'd36105: data <= 8'h00;
            16'd36106: data <= 8'h1F;
            16'd36107: data <= 8'h00;
            16'd36108: data <= 8'h1F;
            16'd36109: data <= 8'h00;
            16'd36110: data <= 8'h1F;
            16'd36111: data <= 8'h00;
            16'd36112: data <= 8'h1F;
            16'd36113: data <= 8'h00;
            16'd36114: data <= 8'h1F;
            16'd36115: data <= 8'h00;
            16'd36116: data <= 8'h1F;
            16'd36117: data <= 8'h00;
            16'd36118: data <= 8'h1F;
            16'd36119: data <= 8'h00;
            16'd36120: data <= 8'hFF;
            16'd36121: data <= 8'hFF;
            16'd36122: data <= 8'h1F;
            16'd36123: data <= 8'h00;
            16'd36124: data <= 8'h1F;
            16'd36125: data <= 8'h00;
            16'd36126: data <= 8'h1F;
            16'd36127: data <= 8'h00;
            16'd36128: data <= 8'h1F;
            16'd36129: data <= 8'h00;
            16'd36130: data <= 8'h1F;
            16'd36131: data <= 8'h00;
            16'd36132: data <= 8'h1F;
            16'd36133: data <= 8'h00;
            16'd36134: data <= 8'h1F;
            16'd36135: data <= 8'h00;
            16'd36136: data <= 8'h1F;
            16'd36137: data <= 8'h00;
            16'd36138: data <= 8'h1F;
            16'd36139: data <= 8'h00;
            16'd36140: data <= 8'h1F;
            16'd36141: data <= 8'h00;
            16'd36142: data <= 8'h1F;
            16'd36143: data <= 8'h00;
            16'd36144: data <= 8'h1F;
            16'd36145: data <= 8'h00;
            16'd36146: data <= 8'h1F;
            16'd36147: data <= 8'h00;
            16'd36148: data <= 8'h1F;
            16'd36149: data <= 8'h00;
            16'd36150: data <= 8'h1F;
            16'd36151: data <= 8'h00;
            16'd36152: data <= 8'h1F;
            16'd36153: data <= 8'h00;
            16'd36154: data <= 8'h1F;
            16'd36155: data <= 8'h00;
            16'd36156: data <= 8'h1F;
            16'd36157: data <= 8'h00;
            16'd36158: data <= 8'h1F;
            16'd36159: data <= 8'h00;
            16'd36160: data <= 8'hFF;
            16'd36161: data <= 8'hFF;
            16'd36162: data <= 8'h1F;
            16'd36163: data <= 8'h00;
            16'd36164: data <= 8'h1F;
            16'd36165: data <= 8'h00;
            16'd36166: data <= 8'h1F;
            16'd36167: data <= 8'h00;
            16'd36168: data <= 8'h1F;
            16'd36169: data <= 8'h00;
            16'd36170: data <= 8'h1F;
            16'd36171: data <= 8'h00;
            16'd36172: data <= 8'h1F;
            16'd36173: data <= 8'h00;
            16'd36174: data <= 8'h1F;
            16'd36175: data <= 8'h00;
            16'd36176: data <= 8'h1F;
            16'd36177: data <= 8'h00;
            16'd36178: data <= 8'h1F;
            16'd36179: data <= 8'h00;
            16'd36180: data <= 8'h1F;
            16'd36181: data <= 8'h00;
            16'd36182: data <= 8'h1F;
            16'd36183: data <= 8'h00;
            16'd36184: data <= 8'h1F;
            16'd36185: data <= 8'h00;
            16'd36186: data <= 8'h1F;
            16'd36187: data <= 8'h00;
            16'd36188: data <= 8'h1F;
            16'd36189: data <= 8'h00;
            16'd36190: data <= 8'h1F;
            16'd36191: data <= 8'h00;
            16'd36192: data <= 8'h1F;
            16'd36193: data <= 8'h00;
            16'd36194: data <= 8'h1F;
            16'd36195: data <= 8'h00;
            16'd36196: data <= 8'h1F;
            16'd36197: data <= 8'h00;
            16'd36198: data <= 8'h1F;
            16'd36199: data <= 8'h00;
            16'd36200: data <= 8'hFF;
            16'd36201: data <= 8'hFF;
            16'd36202: data <= 8'h1F;
            16'd36203: data <= 8'h00;
            16'd36204: data <= 8'h1F;
            16'd36205: data <= 8'h00;
            16'd36206: data <= 8'h1F;
            16'd36207: data <= 8'h00;
            16'd36208: data <= 8'h1F;
            16'd36209: data <= 8'h00;
            16'd36210: data <= 8'h1F;
            16'd36211: data <= 8'h00;
            16'd36212: data <= 8'h1F;
            16'd36213: data <= 8'h00;
            16'd36214: data <= 8'h1F;
            16'd36215: data <= 8'h00;
            16'd36216: data <= 8'h1F;
            16'd36217: data <= 8'h00;
            16'd36218: data <= 8'h1F;
            16'd36219: data <= 8'h00;
            16'd36220: data <= 8'h1F;
            16'd36221: data <= 8'h00;
            16'd36222: data <= 8'h1F;
            16'd36223: data <= 8'h00;
            16'd36224: data <= 8'h1F;
            16'd36225: data <= 8'h00;
            16'd36226: data <= 8'h1F;
            16'd36227: data <= 8'h00;
            16'd36228: data <= 8'h1F;
            16'd36229: data <= 8'h00;
            16'd36230: data <= 8'h1F;
            16'd36231: data <= 8'h00;
            16'd36232: data <= 8'h1F;
            16'd36233: data <= 8'h00;
            16'd36234: data <= 8'h1F;
            16'd36235: data <= 8'h00;
            16'd36236: data <= 8'h1F;
            16'd36237: data <= 8'h00;
            16'd36238: data <= 8'h1F;
            16'd36239: data <= 8'h00;
            16'd36240: data <= 8'hFF;
            16'd36241: data <= 8'hFF;
            16'd36242: data <= 8'h1F;
            16'd36243: data <= 8'h00;
            16'd36244: data <= 8'h1F;
            16'd36245: data <= 8'h00;
            16'd36246: data <= 8'h1F;
            16'd36247: data <= 8'h00;
            16'd36248: data <= 8'h1F;
            16'd36249: data <= 8'h00;
            16'd36250: data <= 8'h1F;
            16'd36251: data <= 8'h00;
            16'd36252: data <= 8'h1F;
            16'd36253: data <= 8'h00;
            16'd36254: data <= 8'h1F;
            16'd36255: data <= 8'h00;
            16'd36256: data <= 8'h1F;
            16'd36257: data <= 8'h00;
            16'd36258: data <= 8'h1F;
            16'd36259: data <= 8'h00;
            16'd36260: data <= 8'h1F;
            16'd36261: data <= 8'h00;
            16'd36262: data <= 8'h1F;
            16'd36263: data <= 8'h00;
            16'd36264: data <= 8'h1F;
            16'd36265: data <= 8'h00;
            16'd36266: data <= 8'h1F;
            16'd36267: data <= 8'h00;
            16'd36268: data <= 8'h1F;
            16'd36269: data <= 8'h00;
            16'd36270: data <= 8'h1F;
            16'd36271: data <= 8'h00;
            16'd36272: data <= 8'h1F;
            16'd36273: data <= 8'h00;
            16'd36274: data <= 8'h1F;
            16'd36275: data <= 8'h00;
            16'd36276: data <= 8'h1F;
            16'd36277: data <= 8'h00;
            16'd36278: data <= 8'h1F;
            16'd36279: data <= 8'h00;
            16'd36280: data <= 8'hFF;
            16'd36281: data <= 8'hFF;
            16'd36282: data <= 8'h1F;
            16'd36283: data <= 8'h00;
            16'd36284: data <= 8'h1F;
            16'd36285: data <= 8'h00;
            16'd36286: data <= 8'h1F;
            16'd36287: data <= 8'h00;
            16'd36288: data <= 8'h1F;
            16'd36289: data <= 8'h00;
            16'd36290: data <= 8'h1F;
            16'd36291: data <= 8'h00;
            16'd36292: data <= 8'h1F;
            16'd36293: data <= 8'h00;
            16'd36294: data <= 8'h1F;
            16'd36295: data <= 8'h00;
            16'd36296: data <= 8'h1F;
            16'd36297: data <= 8'h00;
            16'd36298: data <= 8'h1F;
            16'd36299: data <= 8'h00;
            16'd36300: data <= 8'h1F;
            16'd36301: data <= 8'h00;
            16'd36302: data <= 8'h1F;
            16'd36303: data <= 8'h00;
            16'd36304: data <= 8'h1F;
            16'd36305: data <= 8'h00;
            16'd36306: data <= 8'h1F;
            16'd36307: data <= 8'h00;
            16'd36308: data <= 8'h1F;
            16'd36309: data <= 8'h00;
            16'd36310: data <= 8'h1F;
            16'd36311: data <= 8'h00;
            16'd36312: data <= 8'h1F;
            16'd36313: data <= 8'h00;
            16'd36314: data <= 8'h1F;
            16'd36315: data <= 8'h00;
            16'd36316: data <= 8'h1F;
            16'd36317: data <= 8'h00;
            16'd36318: data <= 8'h1F;
            16'd36319: data <= 8'h00;
            16'd36320: data <= 8'hFF;
            16'd36321: data <= 8'hFF;
            16'd36322: data <= 8'h1F;
            16'd36323: data <= 8'h00;
            16'd36324: data <= 8'h1F;
            16'd36325: data <= 8'h00;
            16'd36326: data <= 8'h1F;
            16'd36327: data <= 8'h00;
            16'd36328: data <= 8'h1F;
            16'd36329: data <= 8'h00;
            16'd36330: data <= 8'h1F;
            16'd36331: data <= 8'h00;
            16'd36332: data <= 8'h1F;
            16'd36333: data <= 8'h00;
            16'd36334: data <= 8'h1F;
            16'd36335: data <= 8'h00;
            16'd36336: data <= 8'h1F;
            16'd36337: data <= 8'h00;
            16'd36338: data <= 8'h1F;
            16'd36339: data <= 8'h00;
            16'd36340: data <= 8'h1F;
            16'd36341: data <= 8'h00;
            16'd36342: data <= 8'h1F;
            16'd36343: data <= 8'h00;
            16'd36344: data <= 8'h1F;
            16'd36345: data <= 8'h00;
            16'd36346: data <= 8'h1F;
            16'd36347: data <= 8'h00;
            16'd36348: data <= 8'h1F;
            16'd36349: data <= 8'h00;
            16'd36350: data <= 8'h1F;
            16'd36351: data <= 8'h00;
            16'd36352: data <= 8'h1F;
            16'd36353: data <= 8'h00;
            16'd36354: data <= 8'h1F;
            16'd36355: data <= 8'h00;
            16'd36356: data <= 8'h1F;
            16'd36357: data <= 8'h00;
            16'd36358: data <= 8'h1F;
            16'd36359: data <= 8'h00;
            16'd36360: data <= 8'hFF;
            16'd36361: data <= 8'hFF;
            16'd36362: data <= 8'h1F;
            16'd36363: data <= 8'h00;
            16'd36364: data <= 8'h1F;
            16'd36365: data <= 8'h00;
            16'd36366: data <= 8'h1F;
            16'd36367: data <= 8'h00;
            16'd36368: data <= 8'h1F;
            16'd36369: data <= 8'h00;
            16'd36370: data <= 8'h1F;
            16'd36371: data <= 8'h00;
            16'd36372: data <= 8'h1F;
            16'd36373: data <= 8'h00;
            16'd36374: data <= 8'h1F;
            16'd36375: data <= 8'h00;
            16'd36376: data <= 8'h1F;
            16'd36377: data <= 8'h00;
            16'd36378: data <= 8'h1F;
            16'd36379: data <= 8'h00;
            16'd36380: data <= 8'h1F;
            16'd36381: data <= 8'h00;
            16'd36382: data <= 8'h1F;
            16'd36383: data <= 8'h00;
            16'd36384: data <= 8'h1F;
            16'd36385: data <= 8'h00;
            16'd36386: data <= 8'h1F;
            16'd36387: data <= 8'h00;
            16'd36388: data <= 8'h1F;
            16'd36389: data <= 8'h00;
            16'd36390: data <= 8'h1F;
            16'd36391: data <= 8'h00;
            16'd36392: data <= 8'h1F;
            16'd36393: data <= 8'h00;
            16'd36394: data <= 8'h1F;
            16'd36395: data <= 8'h00;
            16'd36396: data <= 8'h1F;
            16'd36397: data <= 8'h00;
            16'd36398: data <= 8'h1F;
            16'd36399: data <= 8'h00;
            16'd36400: data <= 8'hFF;
            16'd36401: data <= 8'hFF;
            16'd36402: data <= 8'h1F;
            16'd36403: data <= 8'h00;
            16'd36404: data <= 8'h1F;
            16'd36405: data <= 8'h00;
            16'd36406: data <= 8'h1F;
            16'd36407: data <= 8'h00;
            16'd36408: data <= 8'h1F;
            16'd36409: data <= 8'h00;
            16'd36410: data <= 8'h1F;
            16'd36411: data <= 8'h00;
            16'd36412: data <= 8'h1F;
            16'd36413: data <= 8'h00;
            16'd36414: data <= 8'h1F;
            16'd36415: data <= 8'h00;
            16'd36416: data <= 8'h1F;
            16'd36417: data <= 8'h00;
            16'd36418: data <= 8'h1F;
            16'd36419: data <= 8'h00;
            16'd36420: data <= 8'h1F;
            16'd36421: data <= 8'h00;
            16'd36422: data <= 8'h1F;
            16'd36423: data <= 8'h00;
            16'd36424: data <= 8'h1F;
            16'd36425: data <= 8'h00;
            16'd36426: data <= 8'h1F;
            16'd36427: data <= 8'h00;
            16'd36428: data <= 8'h1F;
            16'd36429: data <= 8'h00;
            16'd36430: data <= 8'h1F;
            16'd36431: data <= 8'h00;
            16'd36432: data <= 8'h1F;
            16'd36433: data <= 8'h00;
            16'd36434: data <= 8'h1F;
            16'd36435: data <= 8'h00;
            16'd36436: data <= 8'h1F;
            16'd36437: data <= 8'h00;
            16'd36438: data <= 8'h1F;
            16'd36439: data <= 8'h00;
            16'd36440: data <= 8'hFF;
            16'd36441: data <= 8'hFF;
            16'd36442: data <= 8'h1F;
            16'd36443: data <= 8'h00;
            16'd36444: data <= 8'h1F;
            16'd36445: data <= 8'h00;
            16'd36446: data <= 8'h1F;
            16'd36447: data <= 8'h00;
            16'd36448: data <= 8'h1F;
            16'd36449: data <= 8'h00;
            16'd36450: data <= 8'h1F;
            16'd36451: data <= 8'h00;
            16'd36452: data <= 8'h1F;
            16'd36453: data <= 8'h00;
            16'd36454: data <= 8'h1F;
            16'd36455: data <= 8'h00;
            16'd36456: data <= 8'h1F;
            16'd36457: data <= 8'h00;
            16'd36458: data <= 8'h1F;
            16'd36459: data <= 8'h00;
            16'd36460: data <= 8'h1F;
            16'd36461: data <= 8'h00;
            16'd36462: data <= 8'h1F;
            16'd36463: data <= 8'h00;
            16'd36464: data <= 8'h1F;
            16'd36465: data <= 8'h00;
            16'd36466: data <= 8'h1F;
            16'd36467: data <= 8'h00;
            16'd36468: data <= 8'h1F;
            16'd36469: data <= 8'h00;
            16'd36470: data <= 8'h1F;
            16'd36471: data <= 8'h00;
            16'd36472: data <= 8'h1F;
            16'd36473: data <= 8'h00;
            16'd36474: data <= 8'h1F;
            16'd36475: data <= 8'h00;
            16'd36476: data <= 8'h1F;
            16'd36477: data <= 8'h00;
            16'd36478: data <= 8'h1F;
            16'd36479: data <= 8'h00;
            16'd36480: data <= 8'hFF;
            16'd36481: data <= 8'hFF;
            16'd36482: data <= 8'h1F;
            16'd36483: data <= 8'h00;
            16'd36484: data <= 8'h1F;
            16'd36485: data <= 8'h00;
            16'd36486: data <= 8'h1F;
            16'd36487: data <= 8'h00;
            16'd36488: data <= 8'h1F;
            16'd36489: data <= 8'h00;
            16'd36490: data <= 8'h1F;
            16'd36491: data <= 8'h00;
            16'd36492: data <= 8'h1F;
            16'd36493: data <= 8'h00;
            16'd36494: data <= 8'h1F;
            16'd36495: data <= 8'h00;
            16'd36496: data <= 8'h1F;
            16'd36497: data <= 8'h00;
            16'd36498: data <= 8'h1F;
            16'd36499: data <= 8'h00;
            16'd36500: data <= 8'h1F;
            16'd36501: data <= 8'h00;
            16'd36502: data <= 8'h1F;
            16'd36503: data <= 8'h00;
            16'd36504: data <= 8'h1F;
            16'd36505: data <= 8'h00;
            16'd36506: data <= 8'h1F;
            16'd36507: data <= 8'h00;
            16'd36508: data <= 8'h1F;
            16'd36509: data <= 8'h00;
            16'd36510: data <= 8'h1F;
            16'd36511: data <= 8'h00;
            16'd36512: data <= 8'h1F;
            16'd36513: data <= 8'h00;
            16'd36514: data <= 8'h1F;
            16'd36515: data <= 8'h00;
            16'd36516: data <= 8'h1F;
            16'd36517: data <= 8'h00;
            16'd36518: data <= 8'h1F;
            16'd36519: data <= 8'h00;
            16'd36520: data <= 8'hFF;
            16'd36521: data <= 8'hFF;
            16'd36522: data <= 8'h1F;
            16'd36523: data <= 8'h00;
            16'd36524: data <= 8'h1F;
            16'd36525: data <= 8'h00;
            16'd36526: data <= 8'h1F;
            16'd36527: data <= 8'h00;
            16'd36528: data <= 8'h1F;
            16'd36529: data <= 8'h00;
            16'd36530: data <= 8'h1F;
            16'd36531: data <= 8'h00;
            16'd36532: data <= 8'h1F;
            16'd36533: data <= 8'h00;
            16'd36534: data <= 8'h1F;
            16'd36535: data <= 8'h00;
            16'd36536: data <= 8'h1F;
            16'd36537: data <= 8'h00;
            16'd36538: data <= 8'h1F;
            16'd36539: data <= 8'h00;
            16'd36540: data <= 8'h1F;
            16'd36541: data <= 8'h00;
            16'd36542: data <= 8'h1F;
            16'd36543: data <= 8'h00;
            16'd36544: data <= 8'h1F;
            16'd36545: data <= 8'h00;
            16'd36546: data <= 8'h1F;
            16'd36547: data <= 8'h00;
            16'd36548: data <= 8'h1F;
            16'd36549: data <= 8'h00;
            16'd36550: data <= 8'h1F;
            16'd36551: data <= 8'h00;
            16'd36552: data <= 8'h1F;
            16'd36553: data <= 8'h00;
            16'd36554: data <= 8'h1F;
            16'd36555: data <= 8'h00;
            16'd36556: data <= 8'h1F;
            16'd36557: data <= 8'h00;
            16'd36558: data <= 8'h1F;
            16'd36559: data <= 8'h00;
            16'd36560: data <= 8'hFF;
            16'd36561: data <= 8'hFF;
            16'd36562: data <= 8'h1F;
            16'd36563: data <= 8'h00;
            16'd36564: data <= 8'h1F;
            16'd36565: data <= 8'h00;
            16'd36566: data <= 8'h1F;
            16'd36567: data <= 8'h00;
            16'd36568: data <= 8'h1F;
            16'd36569: data <= 8'h00;
            16'd36570: data <= 8'h1F;
            16'd36571: data <= 8'h00;
            16'd36572: data <= 8'h1F;
            16'd36573: data <= 8'h00;
            16'd36574: data <= 8'h1F;
            16'd36575: data <= 8'h00;
            16'd36576: data <= 8'h1F;
            16'd36577: data <= 8'h00;
            16'd36578: data <= 8'h1F;
            16'd36579: data <= 8'h00;
            16'd36580: data <= 8'h1F;
            16'd36581: data <= 8'h00;
            16'd36582: data <= 8'h1F;
            16'd36583: data <= 8'h00;
            16'd36584: data <= 8'h1F;
            16'd36585: data <= 8'h00;
            16'd36586: data <= 8'h1F;
            16'd36587: data <= 8'h00;
            16'd36588: data <= 8'h1F;
            16'd36589: data <= 8'h00;
            16'd36590: data <= 8'h1F;
            16'd36591: data <= 8'h00;
            16'd36592: data <= 8'h1F;
            16'd36593: data <= 8'h00;
            16'd36594: data <= 8'h1F;
            16'd36595: data <= 8'h00;
            16'd36596: data <= 8'h1F;
            16'd36597: data <= 8'h00;
            16'd36598: data <= 8'h1F;
            16'd36599: data <= 8'h00;
            16'd36600: data <= 8'hFF;
            16'd36601: data <= 8'hFF;
            16'd36602: data <= 8'h1F;
            16'd36603: data <= 8'h00;
            16'd36604: data <= 8'h1F;
            16'd36605: data <= 8'h00;
            16'd36606: data <= 8'h1F;
            16'd36607: data <= 8'h00;
            16'd36608: data <= 8'h1F;
            16'd36609: data <= 8'h00;
            16'd36610: data <= 8'h1F;
            16'd36611: data <= 8'h00;
            16'd36612: data <= 8'h1F;
            16'd36613: data <= 8'h00;
            16'd36614: data <= 8'h1F;
            16'd36615: data <= 8'h00;
            16'd36616: data <= 8'h1F;
            16'd36617: data <= 8'h00;
            16'd36618: data <= 8'h1F;
            16'd36619: data <= 8'h00;
            16'd36620: data <= 8'h1F;
            16'd36621: data <= 8'h00;
            16'd36622: data <= 8'h1F;
            16'd36623: data <= 8'h00;
            16'd36624: data <= 8'h1F;
            16'd36625: data <= 8'h00;
            16'd36626: data <= 8'h1F;
            16'd36627: data <= 8'h00;
            16'd36628: data <= 8'h1F;
            16'd36629: data <= 8'h00;
            16'd36630: data <= 8'h1F;
            16'd36631: data <= 8'h00;
            16'd36632: data <= 8'h1F;
            16'd36633: data <= 8'h00;
            16'd36634: data <= 8'h1F;
            16'd36635: data <= 8'h00;
            16'd36636: data <= 8'h1F;
            16'd36637: data <= 8'h00;
            16'd36638: data <= 8'h1F;
            16'd36639: data <= 8'h00;
            16'd36640: data <= 8'hFF;
            16'd36641: data <= 8'hFF;
            16'd36642: data <= 8'h1F;
            16'd36643: data <= 8'h00;
            16'd36644: data <= 8'h1F;
            16'd36645: data <= 8'h00;
            16'd36646: data <= 8'h1F;
            16'd36647: data <= 8'h00;
            16'd36648: data <= 8'h1F;
            16'd36649: data <= 8'h00;
            16'd36650: data <= 8'h1F;
            16'd36651: data <= 8'h00;
            16'd36652: data <= 8'h1F;
            16'd36653: data <= 8'h00;
            16'd36654: data <= 8'h1F;
            16'd36655: data <= 8'h00;
            16'd36656: data <= 8'h1F;
            16'd36657: data <= 8'h00;
            16'd36658: data <= 8'h1F;
            16'd36659: data <= 8'h00;
            16'd36660: data <= 8'h1F;
            16'd36661: data <= 8'h00;
            16'd36662: data <= 8'h1F;
            16'd36663: data <= 8'h00;
            16'd36664: data <= 8'h1F;
            16'd36665: data <= 8'h00;
            16'd36666: data <= 8'h1F;
            16'd36667: data <= 8'h00;
            16'd36668: data <= 8'h1F;
            16'd36669: data <= 8'h00;
            16'd36670: data <= 8'h1F;
            16'd36671: data <= 8'h00;
            16'd36672: data <= 8'h1F;
            16'd36673: data <= 8'h00;
            16'd36674: data <= 8'h1F;
            16'd36675: data <= 8'h00;
            16'd36676: data <= 8'h1F;
            16'd36677: data <= 8'h00;
            16'd36678: data <= 8'h1F;
            16'd36679: data <= 8'h00;
            16'd36680: data <= 8'hFF;
            16'd36681: data <= 8'hFF;
            16'd36682: data <= 8'h1F;
            16'd36683: data <= 8'h00;
            16'd36684: data <= 8'h1F;
            16'd36685: data <= 8'h00;
            16'd36686: data <= 8'h1F;
            16'd36687: data <= 8'h00;
            16'd36688: data <= 8'h1F;
            16'd36689: data <= 8'h00;
            16'd36690: data <= 8'h1F;
            16'd36691: data <= 8'h00;
            16'd36692: data <= 8'h1F;
            16'd36693: data <= 8'h00;
            16'd36694: data <= 8'h1F;
            16'd36695: data <= 8'h00;
            16'd36696: data <= 8'h1F;
            16'd36697: data <= 8'h00;
            16'd36698: data <= 8'h1F;
            16'd36699: data <= 8'h00;
            16'd36700: data <= 8'h1F;
            16'd36701: data <= 8'h00;
            16'd36702: data <= 8'h1F;
            16'd36703: data <= 8'h00;
            16'd36704: data <= 8'h1F;
            16'd36705: data <= 8'h00;
            16'd36706: data <= 8'h1F;
            16'd36707: data <= 8'h00;
            16'd36708: data <= 8'h1F;
            16'd36709: data <= 8'h00;
            16'd36710: data <= 8'h1F;
            16'd36711: data <= 8'h00;
            16'd36712: data <= 8'h1F;
            16'd36713: data <= 8'h00;
            16'd36714: data <= 8'h1F;
            16'd36715: data <= 8'h00;
            16'd36716: data <= 8'h1F;
            16'd36717: data <= 8'h00;
            16'd36718: data <= 8'h1F;
            16'd36719: data <= 8'h00;
            16'd36720: data <= 8'hFF;
            16'd36721: data <= 8'hFF;
            16'd36722: data <= 8'h1F;
            16'd36723: data <= 8'h00;
            16'd36724: data <= 8'h1F;
            16'd36725: data <= 8'h00;
            16'd36726: data <= 8'h1F;
            16'd36727: data <= 8'h00;
            16'd36728: data <= 8'h1F;
            16'd36729: data <= 8'h00;
            16'd36730: data <= 8'h1F;
            16'd36731: data <= 8'h00;
            16'd36732: data <= 8'h1F;
            16'd36733: data <= 8'h00;
            16'd36734: data <= 8'h1F;
            16'd36735: data <= 8'h00;
            16'd36736: data <= 8'h1F;
            16'd36737: data <= 8'h00;
            16'd36738: data <= 8'h1F;
            16'd36739: data <= 8'h00;
            16'd36740: data <= 8'h1F;
            16'd36741: data <= 8'h00;
            16'd36742: data <= 8'h1F;
            16'd36743: data <= 8'h00;
            16'd36744: data <= 8'h1F;
            16'd36745: data <= 8'h00;
            16'd36746: data <= 8'h1F;
            16'd36747: data <= 8'h00;
            16'd36748: data <= 8'h1F;
            16'd36749: data <= 8'h00;
            16'd36750: data <= 8'h1F;
            16'd36751: data <= 8'h00;
            16'd36752: data <= 8'h1F;
            16'd36753: data <= 8'h00;
            16'd36754: data <= 8'h1F;
            16'd36755: data <= 8'h00;
            16'd36756: data <= 8'h1F;
            16'd36757: data <= 8'h00;
            16'd36758: data <= 8'h1F;
            16'd36759: data <= 8'h00;
            16'd36760: data <= 8'hFF;
            16'd36761: data <= 8'hFF;
            16'd36762: data <= 8'h1F;
            16'd36763: data <= 8'h00;
            16'd36764: data <= 8'h1F;
            16'd36765: data <= 8'h00;
            16'd36766: data <= 8'h1F;
            16'd36767: data <= 8'h00;
            16'd36768: data <= 8'h1F;
            16'd36769: data <= 8'h00;
            16'd36770: data <= 8'h1F;
            16'd36771: data <= 8'h00;
            16'd36772: data <= 8'h1F;
            16'd36773: data <= 8'h00;
            16'd36774: data <= 8'h1F;
            16'd36775: data <= 8'h00;
            16'd36776: data <= 8'h1F;
            16'd36777: data <= 8'h00;
            16'd36778: data <= 8'h1F;
            16'd36779: data <= 8'h00;
            16'd36780: data <= 8'h1F;
            16'd36781: data <= 8'h00;
            16'd36782: data <= 8'h1F;
            16'd36783: data <= 8'h00;
            16'd36784: data <= 8'h1F;
            16'd36785: data <= 8'h00;
            16'd36786: data <= 8'h1F;
            16'd36787: data <= 8'h00;
            16'd36788: data <= 8'h1F;
            16'd36789: data <= 8'h00;
            16'd36790: data <= 8'h1F;
            16'd36791: data <= 8'h00;
            16'd36792: data <= 8'h1F;
            16'd36793: data <= 8'h00;
            16'd36794: data <= 8'h1F;
            16'd36795: data <= 8'h00;
            16'd36796: data <= 8'h1F;
            16'd36797: data <= 8'h00;
            16'd36798: data <= 8'h1F;
            16'd36799: data <= 8'h00;
            16'd36800: data <= 8'hFF;
            16'd36801: data <= 8'hFF;
            16'd36802: data <= 8'h1F;
            16'd36803: data <= 8'h00;
            16'd36804: data <= 8'h1F;
            16'd36805: data <= 8'h00;
            16'd36806: data <= 8'h1F;
            16'd36807: data <= 8'h00;
            16'd36808: data <= 8'h1F;
            16'd36809: data <= 8'h00;
            16'd36810: data <= 8'h1F;
            16'd36811: data <= 8'h00;
            16'd36812: data <= 8'h1F;
            16'd36813: data <= 8'h00;
            16'd36814: data <= 8'h1F;
            16'd36815: data <= 8'h00;
            16'd36816: data <= 8'h1F;
            16'd36817: data <= 8'h00;
            16'd36818: data <= 8'h1F;
            16'd36819: data <= 8'h00;
            16'd36820: data <= 8'h1F;
            16'd36821: data <= 8'h00;
            16'd36822: data <= 8'h1F;
            16'd36823: data <= 8'h00;
            16'd36824: data <= 8'h1F;
            16'd36825: data <= 8'h00;
            16'd36826: data <= 8'h1F;
            16'd36827: data <= 8'h00;
            16'd36828: data <= 8'h1F;
            16'd36829: data <= 8'h00;
            16'd36830: data <= 8'h1F;
            16'd36831: data <= 8'h00;
            16'd36832: data <= 8'h1F;
            16'd36833: data <= 8'h00;
            16'd36834: data <= 8'h1F;
            16'd36835: data <= 8'h00;
            16'd36836: data <= 8'h1F;
            16'd36837: data <= 8'h00;
            16'd36838: data <= 8'h1F;
            16'd36839: data <= 8'h00;
            16'd36840: data <= 8'hFF;
            16'd36841: data <= 8'hFF;
            16'd36842: data <= 8'h1F;
            16'd36843: data <= 8'h00;
            16'd36844: data <= 8'h1F;
            16'd36845: data <= 8'h00;
            16'd36846: data <= 8'h1F;
            16'd36847: data <= 8'h00;
            16'd36848: data <= 8'h1F;
            16'd36849: data <= 8'h00;
            16'd36850: data <= 8'h1F;
            16'd36851: data <= 8'h00;
            16'd36852: data <= 8'h1F;
            16'd36853: data <= 8'h00;
            16'd36854: data <= 8'h1F;
            16'd36855: data <= 8'h00;
            16'd36856: data <= 8'h1F;
            16'd36857: data <= 8'h00;
            16'd36858: data <= 8'h1F;
            16'd36859: data <= 8'h00;
            16'd36860: data <= 8'h1F;
            16'd36861: data <= 8'h00;
            16'd36862: data <= 8'h1F;
            16'd36863: data <= 8'h00;
            16'd36864: data <= 8'h1F;
            16'd36865: data <= 8'h00;
            16'd36866: data <= 8'h1F;
            16'd36867: data <= 8'h00;
            16'd36868: data <= 8'h1F;
            16'd36869: data <= 8'h00;
            16'd36870: data <= 8'h1F;
            16'd36871: data <= 8'h00;
            16'd36872: data <= 8'h1F;
            16'd36873: data <= 8'h00;
            16'd36874: data <= 8'h1F;
            16'd36875: data <= 8'h00;
            16'd36876: data <= 8'h1F;
            16'd36877: data <= 8'h00;
            16'd36878: data <= 8'h1F;
            16'd36879: data <= 8'h00;
            16'd36880: data <= 8'hFF;
            16'd36881: data <= 8'hFF;
            16'd36882: data <= 8'h1F;
            16'd36883: data <= 8'h00;
            16'd36884: data <= 8'h1F;
            16'd36885: data <= 8'h00;
            16'd36886: data <= 8'h1F;
            16'd36887: data <= 8'h00;
            16'd36888: data <= 8'h1F;
            16'd36889: data <= 8'h00;
            16'd36890: data <= 8'h1F;
            16'd36891: data <= 8'h00;
            16'd36892: data <= 8'h1F;
            16'd36893: data <= 8'h00;
            16'd36894: data <= 8'h1F;
            16'd36895: data <= 8'h00;
            16'd36896: data <= 8'h1F;
            16'd36897: data <= 8'h00;
            16'd36898: data <= 8'h1F;
            16'd36899: data <= 8'h00;
            16'd36900: data <= 8'h1F;
            16'd36901: data <= 8'h00;
            16'd36902: data <= 8'h1F;
            16'd36903: data <= 8'h00;
            16'd36904: data <= 8'h1F;
            16'd36905: data <= 8'h00;
            16'd36906: data <= 8'h1F;
            16'd36907: data <= 8'h00;
            16'd36908: data <= 8'h1F;
            16'd36909: data <= 8'h00;
            16'd36910: data <= 8'h1F;
            16'd36911: data <= 8'h00;
            16'd36912: data <= 8'h1F;
            16'd36913: data <= 8'h00;
            16'd36914: data <= 8'h1F;
            16'd36915: data <= 8'h00;
            16'd36916: data <= 8'h1F;
            16'd36917: data <= 8'h00;
            16'd36918: data <= 8'h1F;
            16'd36919: data <= 8'h00;
            16'd36920: data <= 8'hFF;
            16'd36921: data <= 8'hFF;
            16'd36922: data <= 8'h1F;
            16'd36923: data <= 8'h00;
            16'd36924: data <= 8'h1F;
            16'd36925: data <= 8'h00;
            16'd36926: data <= 8'h1F;
            16'd36927: data <= 8'h00;
            16'd36928: data <= 8'h1F;
            16'd36929: data <= 8'h00;
            16'd36930: data <= 8'h1F;
            16'd36931: data <= 8'h00;
            16'd36932: data <= 8'h1F;
            16'd36933: data <= 8'h00;
            16'd36934: data <= 8'h1F;
            16'd36935: data <= 8'h00;
            16'd36936: data <= 8'h1F;
            16'd36937: data <= 8'h00;
            16'd36938: data <= 8'h1F;
            16'd36939: data <= 8'h00;
            16'd36940: data <= 8'h1F;
            16'd36941: data <= 8'h00;
            16'd36942: data <= 8'h1F;
            16'd36943: data <= 8'h00;
            16'd36944: data <= 8'h1F;
            16'd36945: data <= 8'h00;
            16'd36946: data <= 8'h1F;
            16'd36947: data <= 8'h00;
            16'd36948: data <= 8'h1F;
            16'd36949: data <= 8'h00;
            16'd36950: data <= 8'h1F;
            16'd36951: data <= 8'h00;
            16'd36952: data <= 8'h1F;
            16'd36953: data <= 8'h00;
            16'd36954: data <= 8'h1F;
            16'd36955: data <= 8'h00;
            16'd36956: data <= 8'h1F;
            16'd36957: data <= 8'h00;
            16'd36958: data <= 8'h1F;
            16'd36959: data <= 8'h00;
            16'd36960: data <= 8'hFF;
            16'd36961: data <= 8'hFF;
            16'd36962: data <= 8'h1F;
            16'd36963: data <= 8'h00;
            16'd36964: data <= 8'h1F;
            16'd36965: data <= 8'h00;
            16'd36966: data <= 8'h1F;
            16'd36967: data <= 8'h00;
            16'd36968: data <= 8'h1F;
            16'd36969: data <= 8'h00;
            16'd36970: data <= 8'h1F;
            16'd36971: data <= 8'h00;
            16'd36972: data <= 8'h1F;
            16'd36973: data <= 8'h00;
            16'd36974: data <= 8'h1F;
            16'd36975: data <= 8'h00;
            16'd36976: data <= 8'h1F;
            16'd36977: data <= 8'h00;
            16'd36978: data <= 8'h1F;
            16'd36979: data <= 8'h00;
            16'd36980: data <= 8'h1F;
            16'd36981: data <= 8'h00;
            16'd36982: data <= 8'h1F;
            16'd36983: data <= 8'h00;
            16'd36984: data <= 8'h1F;
            16'd36985: data <= 8'h00;
            16'd36986: data <= 8'h1F;
            16'd36987: data <= 8'h00;
            16'd36988: data <= 8'h1F;
            16'd36989: data <= 8'h00;
            16'd36990: data <= 8'h1F;
            16'd36991: data <= 8'h00;
            16'd36992: data <= 8'h1F;
            16'd36993: data <= 8'h00;
            16'd36994: data <= 8'h1F;
            16'd36995: data <= 8'h00;
            16'd36996: data <= 8'h1F;
            16'd36997: data <= 8'h00;
            16'd36998: data <= 8'h1F;
            16'd36999: data <= 8'h00;
            16'd37000: data <= 8'hFF;
            16'd37001: data <= 8'hFF;
            16'd37002: data <= 8'h1F;
            16'd37003: data <= 8'h00;
            16'd37004: data <= 8'h1F;
            16'd37005: data <= 8'h00;
            16'd37006: data <= 8'h1F;
            16'd37007: data <= 8'h00;
            16'd37008: data <= 8'h1F;
            16'd37009: data <= 8'h00;
            16'd37010: data <= 8'h1F;
            16'd37011: data <= 8'h00;
            16'd37012: data <= 8'h1F;
            16'd37013: data <= 8'h00;
            16'd37014: data <= 8'h1F;
            16'd37015: data <= 8'h00;
            16'd37016: data <= 8'h1F;
            16'd37017: data <= 8'h00;
            16'd37018: data <= 8'h1F;
            16'd37019: data <= 8'h00;
            16'd37020: data <= 8'h1F;
            16'd37021: data <= 8'h00;
            16'd37022: data <= 8'h1F;
            16'd37023: data <= 8'h00;
            16'd37024: data <= 8'h1F;
            16'd37025: data <= 8'h00;
            16'd37026: data <= 8'h1F;
            16'd37027: data <= 8'h00;
            16'd37028: data <= 8'h1F;
            16'd37029: data <= 8'h00;
            16'd37030: data <= 8'h1F;
            16'd37031: data <= 8'h00;
            16'd37032: data <= 8'h1F;
            16'd37033: data <= 8'h00;
            16'd37034: data <= 8'h1F;
            16'd37035: data <= 8'h00;
            16'd37036: data <= 8'h1F;
            16'd37037: data <= 8'h00;
            16'd37038: data <= 8'h1F;
            16'd37039: data <= 8'h00;
            16'd37040: data <= 8'hFF;
            16'd37041: data <= 8'hFF;
            16'd37042: data <= 8'h1F;
            16'd37043: data <= 8'h00;
            16'd37044: data <= 8'h1F;
            16'd37045: data <= 8'h00;
            16'd37046: data <= 8'h1F;
            16'd37047: data <= 8'h00;
            16'd37048: data <= 8'h1F;
            16'd37049: data <= 8'h00;
            16'd37050: data <= 8'h1F;
            16'd37051: data <= 8'h00;
            16'd37052: data <= 8'h1F;
            16'd37053: data <= 8'h00;
            16'd37054: data <= 8'h1F;
            16'd37055: data <= 8'h00;
            16'd37056: data <= 8'h1F;
            16'd37057: data <= 8'h00;
            16'd37058: data <= 8'h1F;
            16'd37059: data <= 8'h00;
            16'd37060: data <= 8'h1F;
            16'd37061: data <= 8'h00;
            16'd37062: data <= 8'h1F;
            16'd37063: data <= 8'h00;
            16'd37064: data <= 8'h1F;
            16'd37065: data <= 8'h00;
            16'd37066: data <= 8'h1F;
            16'd37067: data <= 8'h00;
            16'd37068: data <= 8'h1F;
            16'd37069: data <= 8'h00;
            16'd37070: data <= 8'h1F;
            16'd37071: data <= 8'h00;
            16'd37072: data <= 8'h1F;
            16'd37073: data <= 8'h00;
            16'd37074: data <= 8'h1F;
            16'd37075: data <= 8'h00;
            16'd37076: data <= 8'h1F;
            16'd37077: data <= 8'h00;
            16'd37078: data <= 8'h1F;
            16'd37079: data <= 8'h00;
            16'd37080: data <= 8'hFF;
            16'd37081: data <= 8'hFF;
            16'd37082: data <= 8'h1F;
            16'd37083: data <= 8'h00;
            16'd37084: data <= 8'h1F;
            16'd37085: data <= 8'h00;
            16'd37086: data <= 8'h1F;
            16'd37087: data <= 8'h00;
            16'd37088: data <= 8'h1F;
            16'd37089: data <= 8'h00;
            16'd37090: data <= 8'h1F;
            16'd37091: data <= 8'h00;
            16'd37092: data <= 8'h1F;
            16'd37093: data <= 8'h00;
            16'd37094: data <= 8'h1F;
            16'd37095: data <= 8'h00;
            16'd37096: data <= 8'h1F;
            16'd37097: data <= 8'h00;
            16'd37098: data <= 8'h1F;
            16'd37099: data <= 8'h00;
            16'd37100: data <= 8'h1F;
            16'd37101: data <= 8'h00;
            16'd37102: data <= 8'h1F;
            16'd37103: data <= 8'h00;
            16'd37104: data <= 8'h1F;
            16'd37105: data <= 8'h00;
            16'd37106: data <= 8'h1F;
            16'd37107: data <= 8'h00;
            16'd37108: data <= 8'h1F;
            16'd37109: data <= 8'h00;
            16'd37110: data <= 8'h1F;
            16'd37111: data <= 8'h00;
            16'd37112: data <= 8'h1F;
            16'd37113: data <= 8'h00;
            16'd37114: data <= 8'h1F;
            16'd37115: data <= 8'h00;
            16'd37116: data <= 8'h1F;
            16'd37117: data <= 8'h00;
            16'd37118: data <= 8'h1F;
            16'd37119: data <= 8'h00;
            16'd37120: data <= 8'hFF;
            16'd37121: data <= 8'hFF;
            16'd37122: data <= 8'h1F;
            16'd37123: data <= 8'h00;
            16'd37124: data <= 8'h1F;
            16'd37125: data <= 8'h00;
            16'd37126: data <= 8'h1F;
            16'd37127: data <= 8'h00;
            16'd37128: data <= 8'h1F;
            16'd37129: data <= 8'h00;
            16'd37130: data <= 8'h1F;
            16'd37131: data <= 8'h00;
            16'd37132: data <= 8'h1F;
            16'd37133: data <= 8'h00;
            16'd37134: data <= 8'h1F;
            16'd37135: data <= 8'h00;
            16'd37136: data <= 8'h1F;
            16'd37137: data <= 8'h00;
            16'd37138: data <= 8'h1F;
            16'd37139: data <= 8'h00;
            16'd37140: data <= 8'h1F;
            16'd37141: data <= 8'h00;
            16'd37142: data <= 8'h1F;
            16'd37143: data <= 8'h00;
            16'd37144: data <= 8'h1F;
            16'd37145: data <= 8'h00;
            16'd37146: data <= 8'h1F;
            16'd37147: data <= 8'h00;
            16'd37148: data <= 8'h1F;
            16'd37149: data <= 8'h00;
            16'd37150: data <= 8'h1F;
            16'd37151: data <= 8'h00;
            16'd37152: data <= 8'h1F;
            16'd37153: data <= 8'h00;
            16'd37154: data <= 8'h1F;
            16'd37155: data <= 8'h00;
            16'd37156: data <= 8'h1F;
            16'd37157: data <= 8'h00;
            16'd37158: data <= 8'h1F;
            16'd37159: data <= 8'h00;
            16'd37160: data <= 8'hFF;
            16'd37161: data <= 8'hFF;
            16'd37162: data <= 8'h1F;
            16'd37163: data <= 8'h00;
            16'd37164: data <= 8'h1F;
            16'd37165: data <= 8'h00;
            16'd37166: data <= 8'h1F;
            16'd37167: data <= 8'h00;
            16'd37168: data <= 8'h1F;
            16'd37169: data <= 8'h00;
            16'd37170: data <= 8'h1F;
            16'd37171: data <= 8'h00;
            16'd37172: data <= 8'h1F;
            16'd37173: data <= 8'h00;
            16'd37174: data <= 8'h1F;
            16'd37175: data <= 8'h00;
            16'd37176: data <= 8'h1F;
            16'd37177: data <= 8'h00;
            16'd37178: data <= 8'h1F;
            16'd37179: data <= 8'h00;
            16'd37180: data <= 8'h1F;
            16'd37181: data <= 8'h00;
            16'd37182: data <= 8'h1F;
            16'd37183: data <= 8'h00;
            16'd37184: data <= 8'h1F;
            16'd37185: data <= 8'h00;
            16'd37186: data <= 8'h1F;
            16'd37187: data <= 8'h00;
            16'd37188: data <= 8'h1F;
            16'd37189: data <= 8'h00;
            16'd37190: data <= 8'h1F;
            16'd37191: data <= 8'h00;
            16'd37192: data <= 8'h1F;
            16'd37193: data <= 8'h00;
            16'd37194: data <= 8'h1F;
            16'd37195: data <= 8'h00;
            16'd37196: data <= 8'h1F;
            16'd37197: data <= 8'h00;
            16'd37198: data <= 8'h1F;
            16'd37199: data <= 8'h00;
            16'd37200: data <= 8'hFF;
            16'd37201: data <= 8'hFF;
            16'd37202: data <= 8'h1F;
            16'd37203: data <= 8'h00;
            16'd37204: data <= 8'h1F;
            16'd37205: data <= 8'h00;
            16'd37206: data <= 8'h1F;
            16'd37207: data <= 8'h00;
            16'd37208: data <= 8'h1F;
            16'd37209: data <= 8'h00;
            16'd37210: data <= 8'h1F;
            16'd37211: data <= 8'h00;
            16'd37212: data <= 8'h1F;
            16'd37213: data <= 8'h00;
            16'd37214: data <= 8'h1F;
            16'd37215: data <= 8'h00;
            16'd37216: data <= 8'h1F;
            16'd37217: data <= 8'h00;
            16'd37218: data <= 8'h1F;
            16'd37219: data <= 8'h00;
            16'd37220: data <= 8'h1F;
            16'd37221: data <= 8'h00;
            16'd37222: data <= 8'h1F;
            16'd37223: data <= 8'h00;
            16'd37224: data <= 8'h1F;
            16'd37225: data <= 8'h00;
            16'd37226: data <= 8'h1F;
            16'd37227: data <= 8'h00;
            16'd37228: data <= 8'h1F;
            16'd37229: data <= 8'h00;
            16'd37230: data <= 8'h1F;
            16'd37231: data <= 8'h00;
            16'd37232: data <= 8'h1F;
            16'd37233: data <= 8'h00;
            16'd37234: data <= 8'h1F;
            16'd37235: data <= 8'h00;
            16'd37236: data <= 8'h1F;
            16'd37237: data <= 8'h00;
            16'd37238: data <= 8'h1F;
            16'd37239: data <= 8'h00;
            16'd37240: data <= 8'hFF;
            16'd37241: data <= 8'hFF;
            16'd37242: data <= 8'h1F;
            16'd37243: data <= 8'h00;
            16'd37244: data <= 8'h1F;
            16'd37245: data <= 8'h00;
            16'd37246: data <= 8'h1F;
            16'd37247: data <= 8'h00;
            16'd37248: data <= 8'h1F;
            16'd37249: data <= 8'h00;
            16'd37250: data <= 8'h1F;
            16'd37251: data <= 8'h00;
            16'd37252: data <= 8'h1F;
            16'd37253: data <= 8'h00;
            16'd37254: data <= 8'h1F;
            16'd37255: data <= 8'h00;
            16'd37256: data <= 8'h1F;
            16'd37257: data <= 8'h00;
            16'd37258: data <= 8'h1F;
            16'd37259: data <= 8'h00;
            16'd37260: data <= 8'h1F;
            16'd37261: data <= 8'h00;
            16'd37262: data <= 8'h1F;
            16'd37263: data <= 8'h00;
            16'd37264: data <= 8'h1F;
            16'd37265: data <= 8'h00;
            16'd37266: data <= 8'h1F;
            16'd37267: data <= 8'h00;
            16'd37268: data <= 8'h1F;
            16'd37269: data <= 8'h00;
            16'd37270: data <= 8'h1F;
            16'd37271: data <= 8'h00;
            16'd37272: data <= 8'h1F;
            16'd37273: data <= 8'h00;
            16'd37274: data <= 8'h1F;
            16'd37275: data <= 8'h00;
            16'd37276: data <= 8'h1F;
            16'd37277: data <= 8'h00;
            16'd37278: data <= 8'h1F;
            16'd37279: data <= 8'h00;
            16'd37280: data <= 8'hFF;
            16'd37281: data <= 8'hFF;
            16'd37282: data <= 8'h1F;
            16'd37283: data <= 8'h00;
            16'd37284: data <= 8'h1F;
            16'd37285: data <= 8'h00;
            16'd37286: data <= 8'h1F;
            16'd37287: data <= 8'h00;
            16'd37288: data <= 8'h1F;
            16'd37289: data <= 8'h00;
            16'd37290: data <= 8'h1F;
            16'd37291: data <= 8'h00;
            16'd37292: data <= 8'h1F;
            16'd37293: data <= 8'h00;
            16'd37294: data <= 8'h1F;
            16'd37295: data <= 8'h00;
            16'd37296: data <= 8'h1F;
            16'd37297: data <= 8'h00;
            16'd37298: data <= 8'h1F;
            16'd37299: data <= 8'h00;
            16'd37300: data <= 8'h1F;
            16'd37301: data <= 8'h00;
            16'd37302: data <= 8'h1F;
            16'd37303: data <= 8'h00;
            16'd37304: data <= 8'h1F;
            16'd37305: data <= 8'h00;
            16'd37306: data <= 8'h1F;
            16'd37307: data <= 8'h00;
            16'd37308: data <= 8'h1F;
            16'd37309: data <= 8'h00;
            16'd37310: data <= 8'h1F;
            16'd37311: data <= 8'h00;
            16'd37312: data <= 8'h1F;
            16'd37313: data <= 8'h00;
            16'd37314: data <= 8'h1F;
            16'd37315: data <= 8'h00;
            16'd37316: data <= 8'h1F;
            16'd37317: data <= 8'h00;
            16'd37318: data <= 8'h1F;
            16'd37319: data <= 8'h00;
            16'd37320: data <= 8'hFF;
            16'd37321: data <= 8'hFF;
            16'd37322: data <= 8'h1F;
            16'd37323: data <= 8'h00;
            16'd37324: data <= 8'h1F;
            16'd37325: data <= 8'h00;
            16'd37326: data <= 8'h1F;
            16'd37327: data <= 8'h00;
            16'd37328: data <= 8'h1F;
            16'd37329: data <= 8'h00;
            16'd37330: data <= 8'h1F;
            16'd37331: data <= 8'h00;
            16'd37332: data <= 8'h1F;
            16'd37333: data <= 8'h00;
            16'd37334: data <= 8'h1F;
            16'd37335: data <= 8'h00;
            16'd37336: data <= 8'h1F;
            16'd37337: data <= 8'h00;
            16'd37338: data <= 8'h1F;
            16'd37339: data <= 8'h00;
            16'd37340: data <= 8'h1F;
            16'd37341: data <= 8'h00;
            16'd37342: data <= 8'h1F;
            16'd37343: data <= 8'h00;
            16'd37344: data <= 8'h1F;
            16'd37345: data <= 8'h00;
            16'd37346: data <= 8'h1F;
            16'd37347: data <= 8'h00;
            16'd37348: data <= 8'h1F;
            16'd37349: data <= 8'h00;
            16'd37350: data <= 8'h1F;
            16'd37351: data <= 8'h00;
            16'd37352: data <= 8'h1F;
            16'd37353: data <= 8'h00;
            16'd37354: data <= 8'h1F;
            16'd37355: data <= 8'h00;
            16'd37356: data <= 8'h1F;
            16'd37357: data <= 8'h00;
            16'd37358: data <= 8'h1F;
            16'd37359: data <= 8'h00;
            16'd37360: data <= 8'hFF;
            16'd37361: data <= 8'hFF;
            16'd37362: data <= 8'h1F;
            16'd37363: data <= 8'h00;
            16'd37364: data <= 8'h1F;
            16'd37365: data <= 8'h00;
            16'd37366: data <= 8'h1F;
            16'd37367: data <= 8'h00;
            16'd37368: data <= 8'h1F;
            16'd37369: data <= 8'h00;
            16'd37370: data <= 8'h1F;
            16'd37371: data <= 8'h00;
            16'd37372: data <= 8'h1F;
            16'd37373: data <= 8'h00;
            16'd37374: data <= 8'h1F;
            16'd37375: data <= 8'h00;
            16'd37376: data <= 8'h1F;
            16'd37377: data <= 8'h00;
            16'd37378: data <= 8'h1F;
            16'd37379: data <= 8'h00;
            16'd37380: data <= 8'h1F;
            16'd37381: data <= 8'h00;
            16'd37382: data <= 8'h1F;
            16'd37383: data <= 8'h00;
            16'd37384: data <= 8'h1F;
            16'd37385: data <= 8'h00;
            16'd37386: data <= 8'h1F;
            16'd37387: data <= 8'h00;
            16'd37388: data <= 8'h1F;
            16'd37389: data <= 8'h00;
            16'd37390: data <= 8'h1F;
            16'd37391: data <= 8'h00;
            16'd37392: data <= 8'h1F;
            16'd37393: data <= 8'h00;
            16'd37394: data <= 8'h1F;
            16'd37395: data <= 8'h00;
            16'd37396: data <= 8'h1F;
            16'd37397: data <= 8'h00;
            16'd37398: data <= 8'h1F;
            16'd37399: data <= 8'h00;
            16'd37400: data <= 8'hFF;
            16'd37401: data <= 8'hFF;
            16'd37402: data <= 8'h1F;
            16'd37403: data <= 8'h00;
            16'd37404: data <= 8'h1F;
            16'd37405: data <= 8'h00;
            16'd37406: data <= 8'h1F;
            16'd37407: data <= 8'h00;
            16'd37408: data <= 8'h1F;
            16'd37409: data <= 8'h00;
            16'd37410: data <= 8'h1F;
            16'd37411: data <= 8'h00;
            16'd37412: data <= 8'h1F;
            16'd37413: data <= 8'h00;
            16'd37414: data <= 8'h1F;
            16'd37415: data <= 8'h00;
            16'd37416: data <= 8'h1F;
            16'd37417: data <= 8'h00;
            16'd37418: data <= 8'h1F;
            16'd37419: data <= 8'h00;
            16'd37420: data <= 8'h1F;
            16'd37421: data <= 8'h00;
            16'd37422: data <= 8'h1F;
            16'd37423: data <= 8'h00;
            16'd37424: data <= 8'h1F;
            16'd37425: data <= 8'h00;
            16'd37426: data <= 8'h1F;
            16'd37427: data <= 8'h00;
            16'd37428: data <= 8'h1F;
            16'd37429: data <= 8'h00;
            16'd37430: data <= 8'h1F;
            16'd37431: data <= 8'h00;
            16'd37432: data <= 8'h1F;
            16'd37433: data <= 8'h00;
            16'd37434: data <= 8'h1F;
            16'd37435: data <= 8'h00;
            16'd37436: data <= 8'h1F;
            16'd37437: data <= 8'h00;
            16'd37438: data <= 8'h1F;
            16'd37439: data <= 8'h00;
            16'd37440: data <= 8'hFF;
            16'd37441: data <= 8'hFF;
            16'd37442: data <= 8'h1F;
            16'd37443: data <= 8'h00;
            16'd37444: data <= 8'h1F;
            16'd37445: data <= 8'h00;
            16'd37446: data <= 8'h1F;
            16'd37447: data <= 8'h00;
            16'd37448: data <= 8'h1F;
            16'd37449: data <= 8'h00;
            16'd37450: data <= 8'h1F;
            16'd37451: data <= 8'h00;
            16'd37452: data <= 8'h1F;
            16'd37453: data <= 8'h00;
            16'd37454: data <= 8'h1F;
            16'd37455: data <= 8'h00;
            16'd37456: data <= 8'h1F;
            16'd37457: data <= 8'h00;
            16'd37458: data <= 8'h1F;
            16'd37459: data <= 8'h00;
            16'd37460: data <= 8'h1F;
            16'd37461: data <= 8'h00;
            16'd37462: data <= 8'h1F;
            16'd37463: data <= 8'h00;
            16'd37464: data <= 8'h1F;
            16'd37465: data <= 8'h00;
            16'd37466: data <= 8'h1F;
            16'd37467: data <= 8'h00;
            16'd37468: data <= 8'h1F;
            16'd37469: data <= 8'h00;
            16'd37470: data <= 8'h1F;
            16'd37471: data <= 8'h00;
            16'd37472: data <= 8'h1F;
            16'd37473: data <= 8'h00;
            16'd37474: data <= 8'h1F;
            16'd37475: data <= 8'h00;
            16'd37476: data <= 8'h1F;
            16'd37477: data <= 8'h00;
            16'd37478: data <= 8'h1F;
            16'd37479: data <= 8'h00;
            16'd37480: data <= 8'hFF;
            16'd37481: data <= 8'hFF;
            16'd37482: data <= 8'h1F;
            16'd37483: data <= 8'h00;
            16'd37484: data <= 8'h1F;
            16'd37485: data <= 8'h00;
            16'd37486: data <= 8'h1F;
            16'd37487: data <= 8'h00;
            16'd37488: data <= 8'h1F;
            16'd37489: data <= 8'h00;
            16'd37490: data <= 8'h1F;
            16'd37491: data <= 8'h00;
            16'd37492: data <= 8'h1F;
            16'd37493: data <= 8'h00;
            16'd37494: data <= 8'h1F;
            16'd37495: data <= 8'h00;
            16'd37496: data <= 8'h1F;
            16'd37497: data <= 8'h00;
            16'd37498: data <= 8'h1F;
            16'd37499: data <= 8'h00;
            16'd37500: data <= 8'h1F;
            16'd37501: data <= 8'h00;
            16'd37502: data <= 8'h1F;
            16'd37503: data <= 8'h00;
            16'd37504: data <= 8'h1F;
            16'd37505: data <= 8'h00;
            16'd37506: data <= 8'h1F;
            16'd37507: data <= 8'h00;
            16'd37508: data <= 8'h1F;
            16'd37509: data <= 8'h00;
            16'd37510: data <= 8'h1F;
            16'd37511: data <= 8'h00;
            16'd37512: data <= 8'h1F;
            16'd37513: data <= 8'h00;
            16'd37514: data <= 8'h1F;
            16'd37515: data <= 8'h00;
            16'd37516: data <= 8'h1F;
            16'd37517: data <= 8'h00;
            16'd37518: data <= 8'h1F;
            16'd37519: data <= 8'h00;
            16'd37520: data <= 8'hFF;
            16'd37521: data <= 8'hFF;
            16'd37522: data <= 8'h1F;
            16'd37523: data <= 8'h00;
            16'd37524: data <= 8'h1F;
            16'd37525: data <= 8'h00;
            16'd37526: data <= 8'h1F;
            16'd37527: data <= 8'h00;
            16'd37528: data <= 8'h1F;
            16'd37529: data <= 8'h00;
            16'd37530: data <= 8'h1F;
            16'd37531: data <= 8'h00;
            16'd37532: data <= 8'h1F;
            16'd37533: data <= 8'h00;
            16'd37534: data <= 8'h1F;
            16'd37535: data <= 8'h00;
            16'd37536: data <= 8'h1F;
            16'd37537: data <= 8'h00;
            16'd37538: data <= 8'h1F;
            16'd37539: data <= 8'h00;
            16'd37540: data <= 8'h1F;
            16'd37541: data <= 8'h00;
            16'd37542: data <= 8'h1F;
            16'd37543: data <= 8'h00;
            16'd37544: data <= 8'h1F;
            16'd37545: data <= 8'h00;
            16'd37546: data <= 8'h1F;
            16'd37547: data <= 8'h00;
            16'd37548: data <= 8'h1F;
            16'd37549: data <= 8'h00;
            16'd37550: data <= 8'h1F;
            16'd37551: data <= 8'h00;
            16'd37552: data <= 8'h1F;
            16'd37553: data <= 8'h00;
            16'd37554: data <= 8'h1F;
            16'd37555: data <= 8'h00;
            16'd37556: data <= 8'h1F;
            16'd37557: data <= 8'h00;
            16'd37558: data <= 8'h1F;
            16'd37559: data <= 8'h00;
            16'd37560: data <= 8'hFF;
            16'd37561: data <= 8'hFF;
            16'd37562: data <= 8'h1F;
            16'd37563: data <= 8'h00;
            16'd37564: data <= 8'h1F;
            16'd37565: data <= 8'h00;
            16'd37566: data <= 8'h1F;
            16'd37567: data <= 8'h00;
            16'd37568: data <= 8'h1F;
            16'd37569: data <= 8'h00;
            16'd37570: data <= 8'h1F;
            16'd37571: data <= 8'h00;
            16'd37572: data <= 8'h1F;
            16'd37573: data <= 8'h00;
            16'd37574: data <= 8'h1F;
            16'd37575: data <= 8'h00;
            16'd37576: data <= 8'h1F;
            16'd37577: data <= 8'h00;
            16'd37578: data <= 8'h1F;
            16'd37579: data <= 8'h00;
            16'd37580: data <= 8'h1F;
            16'd37581: data <= 8'h00;
            16'd37582: data <= 8'h1F;
            16'd37583: data <= 8'h00;
            16'd37584: data <= 8'h1F;
            16'd37585: data <= 8'h00;
            16'd37586: data <= 8'h1F;
            16'd37587: data <= 8'h00;
            16'd37588: data <= 8'h1F;
            16'd37589: data <= 8'h00;
            16'd37590: data <= 8'h1F;
            16'd37591: data <= 8'h00;
            16'd37592: data <= 8'h1F;
            16'd37593: data <= 8'h00;
            16'd37594: data <= 8'h1F;
            16'd37595: data <= 8'h00;
            16'd37596: data <= 8'h1F;
            16'd37597: data <= 8'h00;
            16'd37598: data <= 8'h1F;
            16'd37599: data <= 8'h00;
            16'd37600: data <= 8'hFF;
            16'd37601: data <= 8'hFF;
            16'd37602: data <= 8'h1F;
            16'd37603: data <= 8'h00;
            16'd37604: data <= 8'h1F;
            16'd37605: data <= 8'h00;
            16'd37606: data <= 8'h1F;
            16'd37607: data <= 8'h00;
            16'd37608: data <= 8'h1F;
            16'd37609: data <= 8'h00;
            16'd37610: data <= 8'h1F;
            16'd37611: data <= 8'h00;
            16'd37612: data <= 8'h1F;
            16'd37613: data <= 8'h00;
            16'd37614: data <= 8'h1F;
            16'd37615: data <= 8'h00;
            16'd37616: data <= 8'h1F;
            16'd37617: data <= 8'h00;
            16'd37618: data <= 8'h1F;
            16'd37619: data <= 8'h00;
            16'd37620: data <= 8'h1F;
            16'd37621: data <= 8'h00;
            16'd37622: data <= 8'h1F;
            16'd37623: data <= 8'h00;
            16'd37624: data <= 8'h1F;
            16'd37625: data <= 8'h00;
            16'd37626: data <= 8'h1F;
            16'd37627: data <= 8'h00;
            16'd37628: data <= 8'h1F;
            16'd37629: data <= 8'h00;
            16'd37630: data <= 8'h1F;
            16'd37631: data <= 8'h00;
            16'd37632: data <= 8'h1F;
            16'd37633: data <= 8'h00;
            16'd37634: data <= 8'h1F;
            16'd37635: data <= 8'h00;
            16'd37636: data <= 8'h1F;
            16'd37637: data <= 8'h00;
            16'd37638: data <= 8'h1F;
            16'd37639: data <= 8'h00;
            16'd37640: data <= 8'hFF;
            16'd37641: data <= 8'hFF;
            16'd37642: data <= 8'h1F;
            16'd37643: data <= 8'h00;
            16'd37644: data <= 8'h1F;
            16'd37645: data <= 8'h00;
            16'd37646: data <= 8'h1F;
            16'd37647: data <= 8'h00;
            16'd37648: data <= 8'h1F;
            16'd37649: data <= 8'h00;
            16'd37650: data <= 8'h1F;
            16'd37651: data <= 8'h00;
            16'd37652: data <= 8'h1F;
            16'd37653: data <= 8'h00;
            16'd37654: data <= 8'h1F;
            16'd37655: data <= 8'h00;
            16'd37656: data <= 8'h1F;
            16'd37657: data <= 8'h00;
            16'd37658: data <= 8'h1F;
            16'd37659: data <= 8'h00;
            16'd37660: data <= 8'h1F;
            16'd37661: data <= 8'h00;
            16'd37662: data <= 8'h1F;
            16'd37663: data <= 8'h00;
            16'd37664: data <= 8'h1F;
            16'd37665: data <= 8'h00;
            16'd37666: data <= 8'h1F;
            16'd37667: data <= 8'h00;
            16'd37668: data <= 8'h1F;
            16'd37669: data <= 8'h00;
            16'd37670: data <= 8'h1F;
            16'd37671: data <= 8'h00;
            16'd37672: data <= 8'h1F;
            16'd37673: data <= 8'h00;
            16'd37674: data <= 8'h1F;
            16'd37675: data <= 8'h00;
            16'd37676: data <= 8'h1F;
            16'd37677: data <= 8'h00;
            16'd37678: data <= 8'h1F;
            16'd37679: data <= 8'h00;
            16'd37680: data <= 8'hFF;
            16'd37681: data <= 8'hFF;
            16'd37682: data <= 8'h1F;
            16'd37683: data <= 8'h00;
            16'd37684: data <= 8'h1F;
            16'd37685: data <= 8'h00;
            16'd37686: data <= 8'h1F;
            16'd37687: data <= 8'h00;
            16'd37688: data <= 8'h1F;
            16'd37689: data <= 8'h00;
            16'd37690: data <= 8'h1F;
            16'd37691: data <= 8'h00;
            16'd37692: data <= 8'h1F;
            16'd37693: data <= 8'h00;
            16'd37694: data <= 8'h1F;
            16'd37695: data <= 8'h00;
            16'd37696: data <= 8'h1F;
            16'd37697: data <= 8'h00;
            16'd37698: data <= 8'h1F;
            16'd37699: data <= 8'h00;
            16'd37700: data <= 8'h1F;
            16'd37701: data <= 8'h00;
            16'd37702: data <= 8'h1F;
            16'd37703: data <= 8'h00;
            16'd37704: data <= 8'h1F;
            16'd37705: data <= 8'h00;
            16'd37706: data <= 8'h1F;
            16'd37707: data <= 8'h00;
            16'd37708: data <= 8'h1F;
            16'd37709: data <= 8'h00;
            16'd37710: data <= 8'h1F;
            16'd37711: data <= 8'h00;
            16'd37712: data <= 8'h1F;
            16'd37713: data <= 8'h00;
            16'd37714: data <= 8'h1F;
            16'd37715: data <= 8'h00;
            16'd37716: data <= 8'h1F;
            16'd37717: data <= 8'h00;
            16'd37718: data <= 8'h1F;
            16'd37719: data <= 8'h00;
            16'd37720: data <= 8'hFF;
            16'd37721: data <= 8'hFF;
            16'd37722: data <= 8'h1F;
            16'd37723: data <= 8'h00;
            16'd37724: data <= 8'h1F;
            16'd37725: data <= 8'h00;
            16'd37726: data <= 8'h1F;
            16'd37727: data <= 8'h00;
            16'd37728: data <= 8'h1F;
            16'd37729: data <= 8'h00;
            16'd37730: data <= 8'h1F;
            16'd37731: data <= 8'h00;
            16'd37732: data <= 8'h1F;
            16'd37733: data <= 8'h00;
            16'd37734: data <= 8'h1F;
            16'd37735: data <= 8'h00;
            16'd37736: data <= 8'h1F;
            16'd37737: data <= 8'h00;
            16'd37738: data <= 8'h1F;
            16'd37739: data <= 8'h00;
            16'd37740: data <= 8'h1F;
            16'd37741: data <= 8'h00;
            16'd37742: data <= 8'h1F;
            16'd37743: data <= 8'h00;
            16'd37744: data <= 8'h1F;
            16'd37745: data <= 8'h00;
            16'd37746: data <= 8'h1F;
            16'd37747: data <= 8'h00;
            16'd37748: data <= 8'h1F;
            16'd37749: data <= 8'h00;
            16'd37750: data <= 8'h1F;
            16'd37751: data <= 8'h00;
            16'd37752: data <= 8'h1F;
            16'd37753: data <= 8'h00;
            16'd37754: data <= 8'h1F;
            16'd37755: data <= 8'h00;
            16'd37756: data <= 8'h1F;
            16'd37757: data <= 8'h00;
            16'd37758: data <= 8'h1F;
            16'd37759: data <= 8'h00;
            16'd37760: data <= 8'hFF;
            16'd37761: data <= 8'hFF;
            16'd37762: data <= 8'h1F;
            16'd37763: data <= 8'h00;
            16'd37764: data <= 8'h1F;
            16'd37765: data <= 8'h00;
            16'd37766: data <= 8'h1F;
            16'd37767: data <= 8'h00;
            16'd37768: data <= 8'h1F;
            16'd37769: data <= 8'h00;
            16'd37770: data <= 8'h1F;
            16'd37771: data <= 8'h00;
            16'd37772: data <= 8'h1F;
            16'd37773: data <= 8'h00;
            16'd37774: data <= 8'h1F;
            16'd37775: data <= 8'h00;
            16'd37776: data <= 8'h1F;
            16'd37777: data <= 8'h00;
            16'd37778: data <= 8'h1F;
            16'd37779: data <= 8'h00;
            16'd37780: data <= 8'h1F;
            16'd37781: data <= 8'h00;
            16'd37782: data <= 8'h1F;
            16'd37783: data <= 8'h00;
            16'd37784: data <= 8'h1F;
            16'd37785: data <= 8'h00;
            16'd37786: data <= 8'h1F;
            16'd37787: data <= 8'h00;
            16'd37788: data <= 8'h1F;
            16'd37789: data <= 8'h00;
            16'd37790: data <= 8'h1F;
            16'd37791: data <= 8'h00;
            16'd37792: data <= 8'h1F;
            16'd37793: data <= 8'h00;
            16'd37794: data <= 8'h1F;
            16'd37795: data <= 8'h00;
            16'd37796: data <= 8'h1F;
            16'd37797: data <= 8'h00;
            16'd37798: data <= 8'h1F;
            16'd37799: data <= 8'h00;
            16'd37800: data <= 8'hFF;
            16'd37801: data <= 8'hFF;
            16'd37802: data <= 8'h1F;
            16'd37803: data <= 8'h00;
            16'd37804: data <= 8'h1F;
            16'd37805: data <= 8'h00;
            16'd37806: data <= 8'h1F;
            16'd37807: data <= 8'h00;
            16'd37808: data <= 8'h1F;
            16'd37809: data <= 8'h00;
            16'd37810: data <= 8'h1F;
            16'd37811: data <= 8'h00;
            16'd37812: data <= 8'h1F;
            16'd37813: data <= 8'h00;
            16'd37814: data <= 8'h1F;
            16'd37815: data <= 8'h00;
            16'd37816: data <= 8'h1F;
            16'd37817: data <= 8'h00;
            16'd37818: data <= 8'h1F;
            16'd37819: data <= 8'h00;
            16'd37820: data <= 8'h1F;
            16'd37821: data <= 8'h00;
            16'd37822: data <= 8'h1F;
            16'd37823: data <= 8'h00;
            16'd37824: data <= 8'h1F;
            16'd37825: data <= 8'h00;
            16'd37826: data <= 8'h1F;
            16'd37827: data <= 8'h00;
            16'd37828: data <= 8'h1F;
            16'd37829: data <= 8'h00;
            16'd37830: data <= 8'h1F;
            16'd37831: data <= 8'h00;
            16'd37832: data <= 8'h1F;
            16'd37833: data <= 8'h00;
            16'd37834: data <= 8'h1F;
            16'd37835: data <= 8'h00;
            16'd37836: data <= 8'h1F;
            16'd37837: data <= 8'h00;
            16'd37838: data <= 8'h1F;
            16'd37839: data <= 8'h00;
            16'd37840: data <= 8'hFF;
            16'd37841: data <= 8'hFF;
            16'd37842: data <= 8'h1F;
            16'd37843: data <= 8'h00;
            16'd37844: data <= 8'h1F;
            16'd37845: data <= 8'h00;
            16'd37846: data <= 8'h1F;
            16'd37847: data <= 8'h00;
            16'd37848: data <= 8'h1F;
            16'd37849: data <= 8'h00;
            16'd37850: data <= 8'h1F;
            16'd37851: data <= 8'h00;
            16'd37852: data <= 8'h1F;
            16'd37853: data <= 8'h00;
            16'd37854: data <= 8'h1F;
            16'd37855: data <= 8'h00;
            16'd37856: data <= 8'h1F;
            16'd37857: data <= 8'h00;
            16'd37858: data <= 8'h1F;
            16'd37859: data <= 8'h00;
            16'd37860: data <= 8'h1F;
            16'd37861: data <= 8'h00;
            16'd37862: data <= 8'h1F;
            16'd37863: data <= 8'h00;
            16'd37864: data <= 8'h1F;
            16'd37865: data <= 8'h00;
            16'd37866: data <= 8'h1F;
            16'd37867: data <= 8'h00;
            16'd37868: data <= 8'h1F;
            16'd37869: data <= 8'h00;
            16'd37870: data <= 8'h1F;
            16'd37871: data <= 8'h00;
            16'd37872: data <= 8'h1F;
            16'd37873: data <= 8'h00;
            16'd37874: data <= 8'h1F;
            16'd37875: data <= 8'h00;
            16'd37876: data <= 8'h1F;
            16'd37877: data <= 8'h00;
            16'd37878: data <= 8'h1F;
            16'd37879: data <= 8'h00;
            16'd37880: data <= 8'hFF;
            16'd37881: data <= 8'hFF;
            16'd37882: data <= 8'h1F;
            16'd37883: data <= 8'h00;
            16'd37884: data <= 8'h1F;
            16'd37885: data <= 8'h00;
            16'd37886: data <= 8'h1F;
            16'd37887: data <= 8'h00;
            16'd37888: data <= 8'h1F;
            16'd37889: data <= 8'h00;
            16'd37890: data <= 8'h1F;
            16'd37891: data <= 8'h00;
            16'd37892: data <= 8'h1F;
            16'd37893: data <= 8'h00;
            16'd37894: data <= 8'h1F;
            16'd37895: data <= 8'h00;
            16'd37896: data <= 8'h1F;
            16'd37897: data <= 8'h00;
            16'd37898: data <= 8'h1F;
            16'd37899: data <= 8'h00;
            16'd37900: data <= 8'h1F;
            16'd37901: data <= 8'h00;
            16'd37902: data <= 8'h1F;
            16'd37903: data <= 8'h00;
            16'd37904: data <= 8'h1F;
            16'd37905: data <= 8'h00;
            16'd37906: data <= 8'h1F;
            16'd37907: data <= 8'h00;
            16'd37908: data <= 8'h1F;
            16'd37909: data <= 8'h00;
            16'd37910: data <= 8'h1F;
            16'd37911: data <= 8'h00;
            16'd37912: data <= 8'h1F;
            16'd37913: data <= 8'h00;
            16'd37914: data <= 8'h1F;
            16'd37915: data <= 8'h00;
            16'd37916: data <= 8'h1F;
            16'd37917: data <= 8'h00;
            16'd37918: data <= 8'h1F;
            16'd37919: data <= 8'h00;
            16'd37920: data <= 8'hFF;
            16'd37921: data <= 8'hFF;
            16'd37922: data <= 8'h1F;
            16'd37923: data <= 8'h00;
            16'd37924: data <= 8'h1F;
            16'd37925: data <= 8'h00;
            16'd37926: data <= 8'h1F;
            16'd37927: data <= 8'h00;
            16'd37928: data <= 8'h1F;
            16'd37929: data <= 8'h00;
            16'd37930: data <= 8'h1F;
            16'd37931: data <= 8'h00;
            16'd37932: data <= 8'h1F;
            16'd37933: data <= 8'h00;
            16'd37934: data <= 8'h1F;
            16'd37935: data <= 8'h00;
            16'd37936: data <= 8'h1F;
            16'd37937: data <= 8'h00;
            16'd37938: data <= 8'h1F;
            16'd37939: data <= 8'h00;
            16'd37940: data <= 8'h1F;
            16'd37941: data <= 8'h00;
            16'd37942: data <= 8'h1F;
            16'd37943: data <= 8'h00;
            16'd37944: data <= 8'h1F;
            16'd37945: data <= 8'h00;
            16'd37946: data <= 8'h1F;
            16'd37947: data <= 8'h00;
            16'd37948: data <= 8'h1F;
            16'd37949: data <= 8'h00;
            16'd37950: data <= 8'h1F;
            16'd37951: data <= 8'h00;
            16'd37952: data <= 8'h1F;
            16'd37953: data <= 8'h00;
            16'd37954: data <= 8'h1F;
            16'd37955: data <= 8'h00;
            16'd37956: data <= 8'h1F;
            16'd37957: data <= 8'h00;
            16'd37958: data <= 8'h1F;
            16'd37959: data <= 8'h00;
            16'd37960: data <= 8'hFF;
            16'd37961: data <= 8'hFF;
            16'd37962: data <= 8'h1F;
            16'd37963: data <= 8'h00;
            16'd37964: data <= 8'h1F;
            16'd37965: data <= 8'h00;
            16'd37966: data <= 8'h1F;
            16'd37967: data <= 8'h00;
            16'd37968: data <= 8'h1F;
            16'd37969: data <= 8'h00;
            16'd37970: data <= 8'h1F;
            16'd37971: data <= 8'h00;
            16'd37972: data <= 8'h1F;
            16'd37973: data <= 8'h00;
            16'd37974: data <= 8'h1F;
            16'd37975: data <= 8'h00;
            16'd37976: data <= 8'h1F;
            16'd37977: data <= 8'h00;
            16'd37978: data <= 8'h1F;
            16'd37979: data <= 8'h00;
            16'd37980: data <= 8'h1F;
            16'd37981: data <= 8'h00;
            16'd37982: data <= 8'h1F;
            16'd37983: data <= 8'h00;
            16'd37984: data <= 8'h1F;
            16'd37985: data <= 8'h00;
            16'd37986: data <= 8'h1F;
            16'd37987: data <= 8'h00;
            16'd37988: data <= 8'h1F;
            16'd37989: data <= 8'h00;
            16'd37990: data <= 8'h1F;
            16'd37991: data <= 8'h00;
            16'd37992: data <= 8'h1F;
            16'd37993: data <= 8'h00;
            16'd37994: data <= 8'h1F;
            16'd37995: data <= 8'h00;
            16'd37996: data <= 8'h1F;
            16'd37997: data <= 8'h00;
            16'd37998: data <= 8'h1F;
            16'd37999: data <= 8'h00;
            16'd38000: data <= 8'hFF;
            16'd38001: data <= 8'hFF;
            16'd38002: data <= 8'h1F;
            16'd38003: data <= 8'h00;
            16'd38004: data <= 8'h1F;
            16'd38005: data <= 8'h00;
            16'd38006: data <= 8'h1F;
            16'd38007: data <= 8'h00;
            16'd38008: data <= 8'h1F;
            16'd38009: data <= 8'h00;
            16'd38010: data <= 8'h1F;
            16'd38011: data <= 8'h00;
            16'd38012: data <= 8'h1F;
            16'd38013: data <= 8'h00;
            16'd38014: data <= 8'h1F;
            16'd38015: data <= 8'h00;
            16'd38016: data <= 8'h1F;
            16'd38017: data <= 8'h00;
            16'd38018: data <= 8'h1F;
            16'd38019: data <= 8'h00;
            16'd38020: data <= 8'h1F;
            16'd38021: data <= 8'h00;
            16'd38022: data <= 8'h1F;
            16'd38023: data <= 8'h00;
            16'd38024: data <= 8'h1F;
            16'd38025: data <= 8'h00;
            16'd38026: data <= 8'h1F;
            16'd38027: data <= 8'h00;
            16'd38028: data <= 8'h1F;
            16'd38029: data <= 8'h00;
            16'd38030: data <= 8'h1F;
            16'd38031: data <= 8'h00;
            16'd38032: data <= 8'h1F;
            16'd38033: data <= 8'h00;
            16'd38034: data <= 8'h1F;
            16'd38035: data <= 8'h00;
            16'd38036: data <= 8'h1F;
            16'd38037: data <= 8'h00;
            16'd38038: data <= 8'h1F;
            16'd38039: data <= 8'h00;
            16'd38040: data <= 8'hFF;
            16'd38041: data <= 8'hFF;
            16'd38042: data <= 8'h1F;
            16'd38043: data <= 8'h00;
            16'd38044: data <= 8'h1F;
            16'd38045: data <= 8'h00;
            16'd38046: data <= 8'h1F;
            16'd38047: data <= 8'h00;
            16'd38048: data <= 8'h1F;
            16'd38049: data <= 8'h00;
            16'd38050: data <= 8'h1F;
            16'd38051: data <= 8'h00;
            16'd38052: data <= 8'h1F;
            16'd38053: data <= 8'h00;
            16'd38054: data <= 8'h1F;
            16'd38055: data <= 8'h00;
            16'd38056: data <= 8'h1F;
            16'd38057: data <= 8'h00;
            16'd38058: data <= 8'h1F;
            16'd38059: data <= 8'h00;
            16'd38060: data <= 8'h1F;
            16'd38061: data <= 8'h00;
            16'd38062: data <= 8'h1F;
            16'd38063: data <= 8'h00;
            16'd38064: data <= 8'h1F;
            16'd38065: data <= 8'h00;
            16'd38066: data <= 8'h1F;
            16'd38067: data <= 8'h00;
            16'd38068: data <= 8'h1F;
            16'd38069: data <= 8'h00;
            16'd38070: data <= 8'h1F;
            16'd38071: data <= 8'h00;
            16'd38072: data <= 8'h1F;
            16'd38073: data <= 8'h00;
            16'd38074: data <= 8'h1F;
            16'd38075: data <= 8'h00;
            16'd38076: data <= 8'h1F;
            16'd38077: data <= 8'h00;
            16'd38078: data <= 8'h1F;
            16'd38079: data <= 8'h00;
            16'd38080: data <= 8'hFF;
            16'd38081: data <= 8'hFF;
            16'd38082: data <= 8'h1F;
            16'd38083: data <= 8'h00;
            16'd38084: data <= 8'h1F;
            16'd38085: data <= 8'h00;
            16'd38086: data <= 8'h1F;
            16'd38087: data <= 8'h00;
            16'd38088: data <= 8'h1F;
            16'd38089: data <= 8'h00;
            16'd38090: data <= 8'h1F;
            16'd38091: data <= 8'h00;
            16'd38092: data <= 8'h1F;
            16'd38093: data <= 8'h00;
            16'd38094: data <= 8'h1F;
            16'd38095: data <= 8'h00;
            16'd38096: data <= 8'h1F;
            16'd38097: data <= 8'h00;
            16'd38098: data <= 8'h1F;
            16'd38099: data <= 8'h00;
            16'd38100: data <= 8'h1F;
            16'd38101: data <= 8'h00;
            16'd38102: data <= 8'h1F;
            16'd38103: data <= 8'h00;
            16'd38104: data <= 8'h1F;
            16'd38105: data <= 8'h00;
            16'd38106: data <= 8'h1F;
            16'd38107: data <= 8'h00;
            16'd38108: data <= 8'h1F;
            16'd38109: data <= 8'h00;
            16'd38110: data <= 8'h1F;
            16'd38111: data <= 8'h00;
            16'd38112: data <= 8'h1F;
            16'd38113: data <= 8'h00;
            16'd38114: data <= 8'h1F;
            16'd38115: data <= 8'h00;
            16'd38116: data <= 8'h1F;
            16'd38117: data <= 8'h00;
            16'd38118: data <= 8'h1F;
            16'd38119: data <= 8'h00;
            16'd38120: data <= 8'hFF;
            16'd38121: data <= 8'hFF;
            16'd38122: data <= 8'h1F;
            16'd38123: data <= 8'h00;
            16'd38124: data <= 8'h1F;
            16'd38125: data <= 8'h00;
            16'd38126: data <= 8'h1F;
            16'd38127: data <= 8'h00;
            16'd38128: data <= 8'h1F;
            16'd38129: data <= 8'h00;
            16'd38130: data <= 8'h1F;
            16'd38131: data <= 8'h00;
            16'd38132: data <= 8'h1F;
            16'd38133: data <= 8'h00;
            16'd38134: data <= 8'h1F;
            16'd38135: data <= 8'h00;
            16'd38136: data <= 8'h1F;
            16'd38137: data <= 8'h00;
            16'd38138: data <= 8'h1F;
            16'd38139: data <= 8'h00;
            16'd38140: data <= 8'h1F;
            16'd38141: data <= 8'h00;
            16'd38142: data <= 8'h1F;
            16'd38143: data <= 8'h00;
            16'd38144: data <= 8'h1F;
            16'd38145: data <= 8'h00;
            16'd38146: data <= 8'h1F;
            16'd38147: data <= 8'h00;
            16'd38148: data <= 8'h1F;
            16'd38149: data <= 8'h00;
            16'd38150: data <= 8'h1F;
            16'd38151: data <= 8'h00;
            16'd38152: data <= 8'h1F;
            16'd38153: data <= 8'h00;
            16'd38154: data <= 8'h1F;
            16'd38155: data <= 8'h00;
            16'd38156: data <= 8'h1F;
            16'd38157: data <= 8'h00;
            16'd38158: data <= 8'h1F;
            16'd38159: data <= 8'h00;
            16'd38160: data <= 8'hFF;
            16'd38161: data <= 8'hFF;
            16'd38162: data <= 8'h1F;
            16'd38163: data <= 8'h00;
            16'd38164: data <= 8'h1F;
            16'd38165: data <= 8'h00;
            16'd38166: data <= 8'h1F;
            16'd38167: data <= 8'h00;
            16'd38168: data <= 8'h1F;
            16'd38169: data <= 8'h00;
            16'd38170: data <= 8'h1F;
            16'd38171: data <= 8'h00;
            16'd38172: data <= 8'h1F;
            16'd38173: data <= 8'h00;
            16'd38174: data <= 8'h1F;
            16'd38175: data <= 8'h00;
            16'd38176: data <= 8'h1F;
            16'd38177: data <= 8'h00;
            16'd38178: data <= 8'h1F;
            16'd38179: data <= 8'h00;
            16'd38180: data <= 8'h1F;
            16'd38181: data <= 8'h00;
            16'd38182: data <= 8'h1F;
            16'd38183: data <= 8'h00;
            16'd38184: data <= 8'h1F;
            16'd38185: data <= 8'h00;
            16'd38186: data <= 8'h1F;
            16'd38187: data <= 8'h00;
            16'd38188: data <= 8'h1F;
            16'd38189: data <= 8'h00;
            16'd38190: data <= 8'h1F;
            16'd38191: data <= 8'h00;
            16'd38192: data <= 8'h1F;
            16'd38193: data <= 8'h00;
            16'd38194: data <= 8'h1F;
            16'd38195: data <= 8'h00;
            16'd38196: data <= 8'h1F;
            16'd38197: data <= 8'h00;
            16'd38198: data <= 8'h1F;
            16'd38199: data <= 8'h00;
            16'd38200: data <= 8'hFF;
            16'd38201: data <= 8'hFF;
            16'd38202: data <= 8'h1F;
            16'd38203: data <= 8'h00;
            16'd38204: data <= 8'h1F;
            16'd38205: data <= 8'h00;
            16'd38206: data <= 8'h1F;
            16'd38207: data <= 8'h00;
            16'd38208: data <= 8'h1F;
            16'd38209: data <= 8'h00;
            16'd38210: data <= 8'h1F;
            16'd38211: data <= 8'h00;
            16'd38212: data <= 8'h1F;
            16'd38213: data <= 8'h00;
            16'd38214: data <= 8'h1F;
            16'd38215: data <= 8'h00;
            16'd38216: data <= 8'h1F;
            16'd38217: data <= 8'h00;
            16'd38218: data <= 8'h1F;
            16'd38219: data <= 8'h00;
            16'd38220: data <= 8'h1F;
            16'd38221: data <= 8'h00;
            16'd38222: data <= 8'h1F;
            16'd38223: data <= 8'h00;
            16'd38224: data <= 8'h1F;
            16'd38225: data <= 8'h00;
            16'd38226: data <= 8'h1F;
            16'd38227: data <= 8'h00;
            16'd38228: data <= 8'h1F;
            16'd38229: data <= 8'h00;
            16'd38230: data <= 8'h1F;
            16'd38231: data <= 8'h00;
            16'd38232: data <= 8'h1F;
            16'd38233: data <= 8'h00;
            16'd38234: data <= 8'h1F;
            16'd38235: data <= 8'h00;
            16'd38236: data <= 8'h1F;
            16'd38237: data <= 8'h00;
            16'd38238: data <= 8'h1F;
            16'd38239: data <= 8'h00;
            16'd38240: data <= 8'hFF;
            16'd38241: data <= 8'hFF;
            16'd38242: data <= 8'h1F;
            16'd38243: data <= 8'h00;
            16'd38244: data <= 8'h1F;
            16'd38245: data <= 8'h00;
            16'd38246: data <= 8'h1F;
            16'd38247: data <= 8'h00;
            16'd38248: data <= 8'h1F;
            16'd38249: data <= 8'h00;
            16'd38250: data <= 8'h1F;
            16'd38251: data <= 8'h00;
            16'd38252: data <= 8'h1F;
            16'd38253: data <= 8'h00;
            16'd38254: data <= 8'h1F;
            16'd38255: data <= 8'h00;
            16'd38256: data <= 8'h1F;
            16'd38257: data <= 8'h00;
            16'd38258: data <= 8'h1F;
            16'd38259: data <= 8'h00;
            16'd38260: data <= 8'h1F;
            16'd38261: data <= 8'h00;
            16'd38262: data <= 8'h1F;
            16'd38263: data <= 8'h00;
            16'd38264: data <= 8'h1F;
            16'd38265: data <= 8'h00;
            16'd38266: data <= 8'h1F;
            16'd38267: data <= 8'h00;
            16'd38268: data <= 8'h1F;
            16'd38269: data <= 8'h00;
            16'd38270: data <= 8'h1F;
            16'd38271: data <= 8'h00;
            16'd38272: data <= 8'h1F;
            16'd38273: data <= 8'h00;
            16'd38274: data <= 8'h1F;
            16'd38275: data <= 8'h00;
            16'd38276: data <= 8'h1F;
            16'd38277: data <= 8'h00;
            16'd38278: data <= 8'h1F;
            16'd38279: data <= 8'h00;
            16'd38280: data <= 8'hFF;
            16'd38281: data <= 8'hFF;
            16'd38282: data <= 8'h1F;
            16'd38283: data <= 8'h00;
            16'd38284: data <= 8'h1F;
            16'd38285: data <= 8'h00;
            16'd38286: data <= 8'h1F;
            16'd38287: data <= 8'h00;
            16'd38288: data <= 8'h1F;
            16'd38289: data <= 8'h00;
            16'd38290: data <= 8'h1F;
            16'd38291: data <= 8'h00;
            16'd38292: data <= 8'h1F;
            16'd38293: data <= 8'h00;
            16'd38294: data <= 8'h1F;
            16'd38295: data <= 8'h00;
            16'd38296: data <= 8'h1F;
            16'd38297: data <= 8'h00;
            16'd38298: data <= 8'h1F;
            16'd38299: data <= 8'h00;
            16'd38300: data <= 8'h1F;
            16'd38301: data <= 8'h00;
            16'd38302: data <= 8'h1F;
            16'd38303: data <= 8'h00;
            16'd38304: data <= 8'h1F;
            16'd38305: data <= 8'h00;
            16'd38306: data <= 8'h1F;
            16'd38307: data <= 8'h00;
            16'd38308: data <= 8'h1F;
            16'd38309: data <= 8'h00;
            16'd38310: data <= 8'h1F;
            16'd38311: data <= 8'h00;
            16'd38312: data <= 8'h1F;
            16'd38313: data <= 8'h00;
            16'd38314: data <= 8'h1F;
            16'd38315: data <= 8'h00;
            16'd38316: data <= 8'h1F;
            16'd38317: data <= 8'h00;
            16'd38318: data <= 8'h1F;
            16'd38319: data <= 8'h00;
            16'd38320: data <= 8'hFF;
            16'd38321: data <= 8'hFF;
            16'd38322: data <= 8'h1F;
            16'd38323: data <= 8'h00;
            16'd38324: data <= 8'h1F;
            16'd38325: data <= 8'h00;
            16'd38326: data <= 8'h1F;
            16'd38327: data <= 8'h00;
            16'd38328: data <= 8'h1F;
            16'd38329: data <= 8'h00;
            16'd38330: data <= 8'h1F;
            16'd38331: data <= 8'h00;
            16'd38332: data <= 8'h1F;
            16'd38333: data <= 8'h00;
            16'd38334: data <= 8'h1F;
            16'd38335: data <= 8'h00;
            16'd38336: data <= 8'h1F;
            16'd38337: data <= 8'h00;
            16'd38338: data <= 8'h1F;
            16'd38339: data <= 8'h00;
            16'd38340: data <= 8'h1F;
            16'd38341: data <= 8'h00;
            16'd38342: data <= 8'h1F;
            16'd38343: data <= 8'h00;
            16'd38344: data <= 8'h1F;
            16'd38345: data <= 8'h00;
            16'd38346: data <= 8'h1F;
            16'd38347: data <= 8'h00;
            16'd38348: data <= 8'h1F;
            16'd38349: data <= 8'h00;
            16'd38350: data <= 8'h1F;
            16'd38351: data <= 8'h00;
            16'd38352: data <= 8'h1F;
            16'd38353: data <= 8'h00;
            16'd38354: data <= 8'h1F;
            16'd38355: data <= 8'h00;
            16'd38356: data <= 8'h1F;
            16'd38357: data <= 8'h00;
            16'd38358: data <= 8'h1F;
            16'd38359: data <= 8'h00;
            16'd38360: data <= 8'hFF;
            16'd38361: data <= 8'hFF;
            16'd38362: data <= 8'h1F;
            16'd38363: data <= 8'h00;
            16'd38364: data <= 8'h1F;
            16'd38365: data <= 8'h00;
            16'd38366: data <= 8'h1F;
            16'd38367: data <= 8'h00;
            16'd38368: data <= 8'h1F;
            16'd38369: data <= 8'h00;
            16'd38370: data <= 8'h1F;
            16'd38371: data <= 8'h00;
            16'd38372: data <= 8'h1F;
            16'd38373: data <= 8'h00;
            16'd38374: data <= 8'h1F;
            16'd38375: data <= 8'h00;
            16'd38376: data <= 8'h1F;
            16'd38377: data <= 8'h00;
            16'd38378: data <= 8'h1F;
            16'd38379: data <= 8'h00;
            16'd38380: data <= 8'h1F;
            16'd38381: data <= 8'h00;
            16'd38382: data <= 8'h1F;
            16'd38383: data <= 8'h00;
            16'd38384: data <= 8'h1F;
            16'd38385: data <= 8'h00;
            16'd38386: data <= 8'h1F;
            16'd38387: data <= 8'h00;
            16'd38388: data <= 8'h1F;
            16'd38389: data <= 8'h00;
            16'd38390: data <= 8'h1F;
            16'd38391: data <= 8'h00;
            16'd38392: data <= 8'h1F;
            16'd38393: data <= 8'h00;
            16'd38394: data <= 8'h1F;
            16'd38395: data <= 8'h00;
            16'd38396: data <= 8'h1F;
            16'd38397: data <= 8'h00;
            16'd38398: data <= 8'h1F;
            16'd38399: data <= 8'h00;
            default: data <= 8'h00;
        endcase
    end

endmodule
