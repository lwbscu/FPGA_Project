// �Զ����ɵĺϲ�ROMģ��
// ����4��ͼƬ��ÿ��240x180
// ��ɫ��ʽ: �ڰ�(1λ)
// ÿ��ͼƬ: 5400 �ֽ�
// �����ݴ�С: 21600 �ֽ�
// ��ַλ��: 15 λ
// ͼƬ�б�: Angry, Angry, Begging, Begging

module combined_images_240x180_rom (
    input wire clk,
    input wire [14:0] addr,
    output reg [7:0] data
);

    // ͼƬ�����ͳߴ����
    parameter TOTAL_IMAGES = 4;
    parameter BYTES_PER_IMAGE = 5400;
    parameter IMAGE_WIDTH = 240;
    parameter IMAGE_HEIGHT = 180;

    // ROM���ݴ洢
    always @(posedge clk) begin
        case (addr)
            15'd0: data <= 8'h00;
            15'd1: data <= 8'h00;
            15'd2: data <= 8'h00;
            15'd3: data <= 8'h00;
            15'd4: data <= 8'h01;
            15'd5: data <= 8'hFF;
            15'd6: data <= 8'hFF;
            15'd7: data <= 8'hFF;
            15'd8: data <= 8'hFF;
            15'd9: data <= 8'hFF;
            15'd10: data <= 8'hFF;
            15'd11: data <= 8'hFF;
            15'd12: data <= 8'hFF;
            15'd13: data <= 8'hFF;
            15'd14: data <= 8'hFF;
            15'd15: data <= 8'hFF;
            15'd16: data <= 8'hFF;
            15'd17: data <= 8'hFF;
            15'd18: data <= 8'hFF;
            15'd19: data <= 8'hFF;
            15'd20: data <= 8'hFF;
            15'd21: data <= 8'hFF;
            15'd22: data <= 8'hFF;
            15'd23: data <= 8'hFF;
            15'd24: data <= 8'hFF;
            15'd25: data <= 8'h80;
            15'd26: data <= 8'h00;
            15'd27: data <= 8'h00;
            15'd28: data <= 8'h00;
            15'd29: data <= 8'h00;
            15'd30: data <= 8'h00;
            15'd31: data <= 8'h00;
            15'd32: data <= 8'h00;
            15'd33: data <= 8'h00;
            15'd34: data <= 8'h01;
            15'd35: data <= 8'hFF;
            15'd36: data <= 8'hFF;
            15'd37: data <= 8'hFF;
            15'd38: data <= 8'hFF;
            15'd39: data <= 8'hFF;
            15'd40: data <= 8'hFF;
            15'd41: data <= 8'hFF;
            15'd42: data <= 8'hFF;
            15'd43: data <= 8'hFF;
            15'd44: data <= 8'hFF;
            15'd45: data <= 8'hFF;
            15'd46: data <= 8'hFF;
            15'd47: data <= 8'hFF;
            15'd48: data <= 8'hFF;
            15'd49: data <= 8'hFF;
            15'd50: data <= 8'hFF;
            15'd51: data <= 8'hFF;
            15'd52: data <= 8'hFF;
            15'd53: data <= 8'hFF;
            15'd54: data <= 8'hFF;
            15'd55: data <= 8'h80;
            15'd56: data <= 8'h00;
            15'd57: data <= 8'h00;
            15'd58: data <= 8'h00;
            15'd59: data <= 8'h00;
            15'd60: data <= 8'h00;
            15'd61: data <= 8'h00;
            15'd62: data <= 8'h00;
            15'd63: data <= 8'h00;
            15'd64: data <= 8'h01;
            15'd65: data <= 8'hFF;
            15'd66: data <= 8'hFF;
            15'd67: data <= 8'hFF;
            15'd68: data <= 8'hFF;
            15'd69: data <= 8'hFF;
            15'd70: data <= 8'hFF;
            15'd71: data <= 8'hFF;
            15'd72: data <= 8'hFF;
            15'd73: data <= 8'hFF;
            15'd74: data <= 8'hFF;
            15'd75: data <= 8'hFF;
            15'd76: data <= 8'hFF;
            15'd77: data <= 8'hFF;
            15'd78: data <= 8'hFF;
            15'd79: data <= 8'hFF;
            15'd80: data <= 8'hFF;
            15'd81: data <= 8'hFF;
            15'd82: data <= 8'hFF;
            15'd83: data <= 8'hFF;
            15'd84: data <= 8'hFF;
            15'd85: data <= 8'h80;
            15'd86: data <= 8'h00;
            15'd87: data <= 8'h00;
            15'd88: data <= 8'h00;
            15'd89: data <= 8'h00;
            15'd90: data <= 8'h00;
            15'd91: data <= 8'h00;
            15'd92: data <= 8'h00;
            15'd93: data <= 8'h00;
            15'd94: data <= 8'h01;
            15'd95: data <= 8'hFF;
            15'd96: data <= 8'hFF;
            15'd97: data <= 8'hFF;
            15'd98: data <= 8'hFF;
            15'd99: data <= 8'hFF;
            15'd100: data <= 8'hFF;
            15'd101: data <= 8'hFF;
            15'd102: data <= 8'hFF;
            15'd103: data <= 8'hFF;
            15'd104: data <= 8'hFF;
            15'd105: data <= 8'hFF;
            15'd106: data <= 8'hFF;
            15'd107: data <= 8'hFF;
            15'd108: data <= 8'hFF;
            15'd109: data <= 8'hFF;
            15'd110: data <= 8'hFF;
            15'd111: data <= 8'hFF;
            15'd112: data <= 8'hFF;
            15'd113: data <= 8'hFF;
            15'd114: data <= 8'hFF;
            15'd115: data <= 8'h80;
            15'd116: data <= 8'h00;
            15'd117: data <= 8'h00;
            15'd118: data <= 8'h00;
            15'd119: data <= 8'h00;
            15'd120: data <= 8'h00;
            15'd121: data <= 8'h00;
            15'd122: data <= 8'h00;
            15'd123: data <= 8'h00;
            15'd124: data <= 8'h01;
            15'd125: data <= 8'hFF;
            15'd126: data <= 8'hFF;
            15'd127: data <= 8'hFF;
            15'd128: data <= 8'hFF;
            15'd129: data <= 8'hFF;
            15'd130: data <= 8'hFF;
            15'd131: data <= 8'hFF;
            15'd132: data <= 8'hFF;
            15'd133: data <= 8'hFF;
            15'd134: data <= 8'hFF;
            15'd135: data <= 8'hFF;
            15'd136: data <= 8'hFF;
            15'd137: data <= 8'hFF;
            15'd138: data <= 8'hFF;
            15'd139: data <= 8'hFF;
            15'd140: data <= 8'hFF;
            15'd141: data <= 8'hFF;
            15'd142: data <= 8'hFF;
            15'd143: data <= 8'hFF;
            15'd144: data <= 8'hFF;
            15'd145: data <= 8'h80;
            15'd146: data <= 8'h00;
            15'd147: data <= 8'h00;
            15'd148: data <= 8'h00;
            15'd149: data <= 8'h00;
            15'd150: data <= 8'h00;
            15'd151: data <= 8'h00;
            15'd152: data <= 8'h00;
            15'd153: data <= 8'h00;
            15'd154: data <= 8'h01;
            15'd155: data <= 8'hFF;
            15'd156: data <= 8'hFF;
            15'd157: data <= 8'hFF;
            15'd158: data <= 8'hFF;
            15'd159: data <= 8'hFF;
            15'd160: data <= 8'hFF;
            15'd161: data <= 8'hFF;
            15'd162: data <= 8'hFF;
            15'd163: data <= 8'hFF;
            15'd164: data <= 8'hFF;
            15'd165: data <= 8'hFF;
            15'd166: data <= 8'hFF;
            15'd167: data <= 8'hFF;
            15'd168: data <= 8'hFF;
            15'd169: data <= 8'hFF;
            15'd170: data <= 8'hFF;
            15'd171: data <= 8'hFF;
            15'd172: data <= 8'hFF;
            15'd173: data <= 8'hFF;
            15'd174: data <= 8'hFF;
            15'd175: data <= 8'h80;
            15'd176: data <= 8'h00;
            15'd177: data <= 8'h00;
            15'd178: data <= 8'h00;
            15'd179: data <= 8'h00;
            15'd180: data <= 8'h00;
            15'd181: data <= 8'h00;
            15'd182: data <= 8'h00;
            15'd183: data <= 8'h00;
            15'd184: data <= 8'h01;
            15'd185: data <= 8'hFF;
            15'd186: data <= 8'hFF;
            15'd187: data <= 8'hFF;
            15'd188: data <= 8'hFF;
            15'd189: data <= 8'hFF;
            15'd190: data <= 8'hFF;
            15'd191: data <= 8'hFF;
            15'd192: data <= 8'hFF;
            15'd193: data <= 8'hFF;
            15'd194: data <= 8'hFF;
            15'd195: data <= 8'hFF;
            15'd196: data <= 8'hFF;
            15'd197: data <= 8'hFF;
            15'd198: data <= 8'hFF;
            15'd199: data <= 8'hFF;
            15'd200: data <= 8'hFF;
            15'd201: data <= 8'hFF;
            15'd202: data <= 8'hFF;
            15'd203: data <= 8'hFF;
            15'd204: data <= 8'hFF;
            15'd205: data <= 8'h80;
            15'd206: data <= 8'h00;
            15'd207: data <= 8'h00;
            15'd208: data <= 8'h00;
            15'd209: data <= 8'h00;
            15'd210: data <= 8'h00;
            15'd211: data <= 8'h00;
            15'd212: data <= 8'h00;
            15'd213: data <= 8'h00;
            15'd214: data <= 8'h01;
            15'd215: data <= 8'hFF;
            15'd216: data <= 8'hFF;
            15'd217: data <= 8'hFF;
            15'd218: data <= 8'hFF;
            15'd219: data <= 8'hFF;
            15'd220: data <= 8'hFF;
            15'd221: data <= 8'hFF;
            15'd222: data <= 8'hFF;
            15'd223: data <= 8'hFF;
            15'd224: data <= 8'hFF;
            15'd225: data <= 8'hFF;
            15'd226: data <= 8'hFF;
            15'd227: data <= 8'hFF;
            15'd228: data <= 8'hFF;
            15'd229: data <= 8'hFF;
            15'd230: data <= 8'hFF;
            15'd231: data <= 8'hFF;
            15'd232: data <= 8'hFF;
            15'd233: data <= 8'hFF;
            15'd234: data <= 8'hFF;
            15'd235: data <= 8'h80;
            15'd236: data <= 8'h00;
            15'd237: data <= 8'h00;
            15'd238: data <= 8'h00;
            15'd239: data <= 8'h00;
            15'd240: data <= 8'h00;
            15'd241: data <= 8'h00;
            15'd242: data <= 8'h00;
            15'd243: data <= 8'h00;
            15'd244: data <= 8'h01;
            15'd245: data <= 8'hFF;
            15'd246: data <= 8'hFF;
            15'd247: data <= 8'hFF;
            15'd248: data <= 8'hFF;
            15'd249: data <= 8'hFF;
            15'd250: data <= 8'hFF;
            15'd251: data <= 8'hFF;
            15'd252: data <= 8'hFF;
            15'd253: data <= 8'hFF;
            15'd254: data <= 8'hFF;
            15'd255: data <= 8'hFF;
            15'd256: data <= 8'hFF;
            15'd257: data <= 8'hFF;
            15'd258: data <= 8'hFF;
            15'd259: data <= 8'hFF;
            15'd260: data <= 8'hFF;
            15'd261: data <= 8'hFF;
            15'd262: data <= 8'hFF;
            15'd263: data <= 8'hFF;
            15'd264: data <= 8'hFF;
            15'd265: data <= 8'h80;
            15'd266: data <= 8'h00;
            15'd267: data <= 8'h00;
            15'd268: data <= 8'h00;
            15'd269: data <= 8'h00;
            15'd270: data <= 8'h00;
            15'd271: data <= 8'h00;
            15'd272: data <= 8'h00;
            15'd273: data <= 8'h00;
            15'd274: data <= 8'h01;
            15'd275: data <= 8'hFF;
            15'd276: data <= 8'hFF;
            15'd277: data <= 8'hFF;
            15'd278: data <= 8'hFF;
            15'd279: data <= 8'hFF;
            15'd280: data <= 8'hFF;
            15'd281: data <= 8'hFF;
            15'd282: data <= 8'hFF;
            15'd283: data <= 8'hFF;
            15'd284: data <= 8'hFF;
            15'd285: data <= 8'hFF;
            15'd286: data <= 8'hFF;
            15'd287: data <= 8'hFF;
            15'd288: data <= 8'hFF;
            15'd289: data <= 8'hFF;
            15'd290: data <= 8'hFF;
            15'd291: data <= 8'hFF;
            15'd292: data <= 8'hFF;
            15'd293: data <= 8'hFF;
            15'd294: data <= 8'hFF;
            15'd295: data <= 8'h80;
            15'd296: data <= 8'h00;
            15'd297: data <= 8'h00;
            15'd298: data <= 8'h00;
            15'd299: data <= 8'h00;
            15'd300: data <= 8'h00;
            15'd301: data <= 8'h00;
            15'd302: data <= 8'h00;
            15'd303: data <= 8'h00;
            15'd304: data <= 8'h01;
            15'd305: data <= 8'hFF;
            15'd306: data <= 8'hFF;
            15'd307: data <= 8'hFF;
            15'd308: data <= 8'hFF;
            15'd309: data <= 8'hFF;
            15'd310: data <= 8'hFF;
            15'd311: data <= 8'hFF;
            15'd312: data <= 8'hFF;
            15'd313: data <= 8'hFF;
            15'd314: data <= 8'hFF;
            15'd315: data <= 8'hFF;
            15'd316: data <= 8'hFF;
            15'd317: data <= 8'hFF;
            15'd318: data <= 8'hFF;
            15'd319: data <= 8'hFF;
            15'd320: data <= 8'hFF;
            15'd321: data <= 8'hFF;
            15'd322: data <= 8'hFF;
            15'd323: data <= 8'hFF;
            15'd324: data <= 8'hFF;
            15'd325: data <= 8'h80;
            15'd326: data <= 8'h00;
            15'd327: data <= 8'h00;
            15'd328: data <= 8'h00;
            15'd329: data <= 8'h00;
            15'd330: data <= 8'h00;
            15'd331: data <= 8'h00;
            15'd332: data <= 8'h00;
            15'd333: data <= 8'h00;
            15'd334: data <= 8'h01;
            15'd335: data <= 8'hFF;
            15'd336: data <= 8'hFF;
            15'd337: data <= 8'hFF;
            15'd338: data <= 8'hFF;
            15'd339: data <= 8'hFF;
            15'd340: data <= 8'hFF;
            15'd341: data <= 8'hFF;
            15'd342: data <= 8'hFF;
            15'd343: data <= 8'hFF;
            15'd344: data <= 8'hFF;
            15'd345: data <= 8'hFF;
            15'd346: data <= 8'hFF;
            15'd347: data <= 8'hFF;
            15'd348: data <= 8'hFF;
            15'd349: data <= 8'hFF;
            15'd350: data <= 8'hFF;
            15'd351: data <= 8'hFF;
            15'd352: data <= 8'hFF;
            15'd353: data <= 8'hFF;
            15'd354: data <= 8'hFF;
            15'd355: data <= 8'h80;
            15'd356: data <= 8'h00;
            15'd357: data <= 8'h00;
            15'd358: data <= 8'h00;
            15'd359: data <= 8'h00;
            15'd360: data <= 8'h00;
            15'd361: data <= 8'h00;
            15'd362: data <= 8'h00;
            15'd363: data <= 8'h00;
            15'd364: data <= 8'h01;
            15'd365: data <= 8'hFF;
            15'd366: data <= 8'hFF;
            15'd367: data <= 8'hFF;
            15'd368: data <= 8'hFF;
            15'd369: data <= 8'hFF;
            15'd370: data <= 8'hFF;
            15'd371: data <= 8'hFF;
            15'd372: data <= 8'hFF;
            15'd373: data <= 8'hFF;
            15'd374: data <= 8'hFF;
            15'd375: data <= 8'hFF;
            15'd376: data <= 8'hFF;
            15'd377: data <= 8'hFF;
            15'd378: data <= 8'hFF;
            15'd379: data <= 8'hFF;
            15'd380: data <= 8'hFF;
            15'd381: data <= 8'hFF;
            15'd382: data <= 8'hFF;
            15'd383: data <= 8'hFF;
            15'd384: data <= 8'hFF;
            15'd385: data <= 8'h80;
            15'd386: data <= 8'h00;
            15'd387: data <= 8'h00;
            15'd388: data <= 8'h00;
            15'd389: data <= 8'h00;
            15'd390: data <= 8'h00;
            15'd391: data <= 8'h00;
            15'd392: data <= 8'h00;
            15'd393: data <= 8'h00;
            15'd394: data <= 8'h01;
            15'd395: data <= 8'hFF;
            15'd396: data <= 8'hFF;
            15'd397: data <= 8'hFF;
            15'd398: data <= 8'hFF;
            15'd399: data <= 8'hFF;
            15'd400: data <= 8'hFF;
            15'd401: data <= 8'hFF;
            15'd402: data <= 8'hFF;
            15'd403: data <= 8'hFF;
            15'd404: data <= 8'hFF;
            15'd405: data <= 8'hFF;
            15'd406: data <= 8'hFF;
            15'd407: data <= 8'hFF;
            15'd408: data <= 8'hFF;
            15'd409: data <= 8'hFF;
            15'd410: data <= 8'hFF;
            15'd411: data <= 8'hFF;
            15'd412: data <= 8'hFF;
            15'd413: data <= 8'hFF;
            15'd414: data <= 8'hFF;
            15'd415: data <= 8'h80;
            15'd416: data <= 8'h00;
            15'd417: data <= 8'h00;
            15'd418: data <= 8'h00;
            15'd419: data <= 8'h00;
            15'd420: data <= 8'h00;
            15'd421: data <= 8'h00;
            15'd422: data <= 8'h00;
            15'd423: data <= 8'h00;
            15'd424: data <= 8'h01;
            15'd425: data <= 8'hFF;
            15'd426: data <= 8'hFF;
            15'd427: data <= 8'hFF;
            15'd428: data <= 8'hFF;
            15'd429: data <= 8'hFF;
            15'd430: data <= 8'hFF;
            15'd431: data <= 8'hFF;
            15'd432: data <= 8'hFF;
            15'd433: data <= 8'hFF;
            15'd434: data <= 8'hFF;
            15'd435: data <= 8'hFF;
            15'd436: data <= 8'hFF;
            15'd437: data <= 8'hFF;
            15'd438: data <= 8'hFF;
            15'd439: data <= 8'hFF;
            15'd440: data <= 8'hFF;
            15'd441: data <= 8'hFF;
            15'd442: data <= 8'hFF;
            15'd443: data <= 8'hFF;
            15'd444: data <= 8'hFF;
            15'd445: data <= 8'h80;
            15'd446: data <= 8'h00;
            15'd447: data <= 8'h00;
            15'd448: data <= 8'h00;
            15'd449: data <= 8'h00;
            15'd450: data <= 8'h00;
            15'd451: data <= 8'h00;
            15'd452: data <= 8'h00;
            15'd453: data <= 8'h00;
            15'd454: data <= 8'h01;
            15'd455: data <= 8'hFF;
            15'd456: data <= 8'hFF;
            15'd457: data <= 8'hFF;
            15'd458: data <= 8'hFF;
            15'd459: data <= 8'hFF;
            15'd460: data <= 8'hFF;
            15'd461: data <= 8'hFF;
            15'd462: data <= 8'hFF;
            15'd463: data <= 8'hFF;
            15'd464: data <= 8'hFF;
            15'd465: data <= 8'hFF;
            15'd466: data <= 8'hFF;
            15'd467: data <= 8'hFF;
            15'd468: data <= 8'hFF;
            15'd469: data <= 8'hFF;
            15'd470: data <= 8'hFF;
            15'd471: data <= 8'hFF;
            15'd472: data <= 8'hFF;
            15'd473: data <= 8'hFF;
            15'd474: data <= 8'hFF;
            15'd475: data <= 8'h80;
            15'd476: data <= 8'h00;
            15'd477: data <= 8'h00;
            15'd478: data <= 8'h00;
            15'd479: data <= 8'h00;
            15'd480: data <= 8'h00;
            15'd481: data <= 8'h00;
            15'd482: data <= 8'h00;
            15'd483: data <= 8'h00;
            15'd484: data <= 8'h01;
            15'd485: data <= 8'hFF;
            15'd486: data <= 8'hFF;
            15'd487: data <= 8'hFF;
            15'd488: data <= 8'hFF;
            15'd489: data <= 8'hFF;
            15'd490: data <= 8'hFF;
            15'd491: data <= 8'hFF;
            15'd492: data <= 8'hFF;
            15'd493: data <= 8'hFF;
            15'd494: data <= 8'hFF;
            15'd495: data <= 8'hFF;
            15'd496: data <= 8'hFF;
            15'd497: data <= 8'hFF;
            15'd498: data <= 8'hFF;
            15'd499: data <= 8'hFF;
            15'd500: data <= 8'hFF;
            15'd501: data <= 8'hFF;
            15'd502: data <= 8'hFF;
            15'd503: data <= 8'hFF;
            15'd504: data <= 8'hFF;
            15'd505: data <= 8'h80;
            15'd506: data <= 8'h00;
            15'd507: data <= 8'h00;
            15'd508: data <= 8'h00;
            15'd509: data <= 8'h00;
            15'd510: data <= 8'h00;
            15'd511: data <= 8'h00;
            15'd512: data <= 8'h00;
            15'd513: data <= 8'h00;
            15'd514: data <= 8'h01;
            15'd515: data <= 8'hFF;
            15'd516: data <= 8'hFF;
            15'd517: data <= 8'hFF;
            15'd518: data <= 8'hFF;
            15'd519: data <= 8'hFF;
            15'd520: data <= 8'hFF;
            15'd521: data <= 8'hFF;
            15'd522: data <= 8'hFF;
            15'd523: data <= 8'hFF;
            15'd524: data <= 8'hFF;
            15'd525: data <= 8'hFF;
            15'd526: data <= 8'hFF;
            15'd527: data <= 8'hFF;
            15'd528: data <= 8'hFF;
            15'd529: data <= 8'hFF;
            15'd530: data <= 8'hFF;
            15'd531: data <= 8'hFF;
            15'd532: data <= 8'hFF;
            15'd533: data <= 8'hFF;
            15'd534: data <= 8'hFF;
            15'd535: data <= 8'h80;
            15'd536: data <= 8'h00;
            15'd537: data <= 8'h00;
            15'd538: data <= 8'h00;
            15'd539: data <= 8'h00;
            15'd540: data <= 8'h00;
            15'd541: data <= 8'h00;
            15'd542: data <= 8'h00;
            15'd543: data <= 8'h00;
            15'd544: data <= 8'h01;
            15'd545: data <= 8'hFF;
            15'd546: data <= 8'hFF;
            15'd547: data <= 8'hFF;
            15'd548: data <= 8'hFF;
            15'd549: data <= 8'hFF;
            15'd550: data <= 8'hFF;
            15'd551: data <= 8'hFF;
            15'd552: data <= 8'hFF;
            15'd553: data <= 8'hFF;
            15'd554: data <= 8'hFF;
            15'd555: data <= 8'hFF;
            15'd556: data <= 8'hFF;
            15'd557: data <= 8'hFF;
            15'd558: data <= 8'hFF;
            15'd559: data <= 8'hFF;
            15'd560: data <= 8'hFF;
            15'd561: data <= 8'hFF;
            15'd562: data <= 8'hFF;
            15'd563: data <= 8'hFF;
            15'd564: data <= 8'hFF;
            15'd565: data <= 8'h80;
            15'd566: data <= 8'h00;
            15'd567: data <= 8'h00;
            15'd568: data <= 8'h00;
            15'd569: data <= 8'h00;
            15'd570: data <= 8'h00;
            15'd571: data <= 8'h00;
            15'd572: data <= 8'h00;
            15'd573: data <= 8'h00;
            15'd574: data <= 8'h01;
            15'd575: data <= 8'hFF;
            15'd576: data <= 8'hFF;
            15'd577: data <= 8'hFF;
            15'd578: data <= 8'hFF;
            15'd579: data <= 8'hFF;
            15'd580: data <= 8'hFF;
            15'd581: data <= 8'hFF;
            15'd582: data <= 8'hFF;
            15'd583: data <= 8'hFF;
            15'd584: data <= 8'hFF;
            15'd585: data <= 8'hFF;
            15'd586: data <= 8'hFF;
            15'd587: data <= 8'hFF;
            15'd588: data <= 8'hFF;
            15'd589: data <= 8'hFF;
            15'd590: data <= 8'hFF;
            15'd591: data <= 8'hFF;
            15'd592: data <= 8'hFF;
            15'd593: data <= 8'hFF;
            15'd594: data <= 8'hFF;
            15'd595: data <= 8'h80;
            15'd596: data <= 8'h00;
            15'd597: data <= 8'h00;
            15'd598: data <= 8'h00;
            15'd599: data <= 8'h00;
            15'd600: data <= 8'h00;
            15'd601: data <= 8'h00;
            15'd602: data <= 8'h00;
            15'd603: data <= 8'h00;
            15'd604: data <= 8'h01;
            15'd605: data <= 8'hFF;
            15'd606: data <= 8'hFF;
            15'd607: data <= 8'hFF;
            15'd608: data <= 8'hFF;
            15'd609: data <= 8'hFF;
            15'd610: data <= 8'hFF;
            15'd611: data <= 8'hFF;
            15'd612: data <= 8'hFF;
            15'd613: data <= 8'hFF;
            15'd614: data <= 8'hFF;
            15'd615: data <= 8'hFF;
            15'd616: data <= 8'hFF;
            15'd617: data <= 8'hFF;
            15'd618: data <= 8'hFF;
            15'd619: data <= 8'hFF;
            15'd620: data <= 8'hFF;
            15'd621: data <= 8'hFF;
            15'd622: data <= 8'hFF;
            15'd623: data <= 8'hFF;
            15'd624: data <= 8'hFF;
            15'd625: data <= 8'h80;
            15'd626: data <= 8'h00;
            15'd627: data <= 8'h00;
            15'd628: data <= 8'h00;
            15'd629: data <= 8'h00;
            15'd630: data <= 8'h00;
            15'd631: data <= 8'h00;
            15'd632: data <= 8'h00;
            15'd633: data <= 8'h00;
            15'd634: data <= 8'h01;
            15'd635: data <= 8'hFF;
            15'd636: data <= 8'hFF;
            15'd637: data <= 8'hFF;
            15'd638: data <= 8'hFF;
            15'd639: data <= 8'hFF;
            15'd640: data <= 8'hFF;
            15'd641: data <= 8'hFF;
            15'd642: data <= 8'hFF;
            15'd643: data <= 8'hFF;
            15'd644: data <= 8'hFF;
            15'd645: data <= 8'hFF;
            15'd646: data <= 8'hFF;
            15'd647: data <= 8'hFF;
            15'd648: data <= 8'hFF;
            15'd649: data <= 8'hFF;
            15'd650: data <= 8'hFF;
            15'd651: data <= 8'hFF;
            15'd652: data <= 8'hFF;
            15'd653: data <= 8'hFF;
            15'd654: data <= 8'hFF;
            15'd655: data <= 8'h80;
            15'd656: data <= 8'h00;
            15'd657: data <= 8'h00;
            15'd658: data <= 8'h00;
            15'd659: data <= 8'h00;
            15'd660: data <= 8'h00;
            15'd661: data <= 8'h00;
            15'd662: data <= 8'h00;
            15'd663: data <= 8'h00;
            15'd664: data <= 8'h01;
            15'd665: data <= 8'hFF;
            15'd666: data <= 8'hFF;
            15'd667: data <= 8'hFF;
            15'd668: data <= 8'hFF;
            15'd669: data <= 8'hFF;
            15'd670: data <= 8'hFF;
            15'd671: data <= 8'hFF;
            15'd672: data <= 8'hFF;
            15'd673: data <= 8'hFF;
            15'd674: data <= 8'hFF;
            15'd675: data <= 8'hFF;
            15'd676: data <= 8'hFF;
            15'd677: data <= 8'hFF;
            15'd678: data <= 8'hFF;
            15'd679: data <= 8'hFF;
            15'd680: data <= 8'hFF;
            15'd681: data <= 8'hFF;
            15'd682: data <= 8'hFF;
            15'd683: data <= 8'hFF;
            15'd684: data <= 8'hFF;
            15'd685: data <= 8'h80;
            15'd686: data <= 8'h00;
            15'd687: data <= 8'h00;
            15'd688: data <= 8'h00;
            15'd689: data <= 8'h00;
            15'd690: data <= 8'h00;
            15'd691: data <= 8'h00;
            15'd692: data <= 8'h00;
            15'd693: data <= 8'h00;
            15'd694: data <= 8'h01;
            15'd695: data <= 8'hFF;
            15'd696: data <= 8'hFF;
            15'd697: data <= 8'hFF;
            15'd698: data <= 8'hFF;
            15'd699: data <= 8'hFF;
            15'd700: data <= 8'hFF;
            15'd701: data <= 8'hFF;
            15'd702: data <= 8'hFF;
            15'd703: data <= 8'hFF;
            15'd704: data <= 8'hFF;
            15'd705: data <= 8'hFF;
            15'd706: data <= 8'hFF;
            15'd707: data <= 8'hFF;
            15'd708: data <= 8'hFF;
            15'd709: data <= 8'hFF;
            15'd710: data <= 8'hFF;
            15'd711: data <= 8'hFF;
            15'd712: data <= 8'hFF;
            15'd713: data <= 8'hFF;
            15'd714: data <= 8'hFF;
            15'd715: data <= 8'h80;
            15'd716: data <= 8'h00;
            15'd717: data <= 8'h00;
            15'd718: data <= 8'h00;
            15'd719: data <= 8'h00;
            15'd720: data <= 8'h00;
            15'd721: data <= 8'h00;
            15'd722: data <= 8'h00;
            15'd723: data <= 8'h00;
            15'd724: data <= 8'h01;
            15'd725: data <= 8'hFF;
            15'd726: data <= 8'hFF;
            15'd727: data <= 8'hFF;
            15'd728: data <= 8'hFF;
            15'd729: data <= 8'hFF;
            15'd730: data <= 8'hFF;
            15'd731: data <= 8'hFF;
            15'd732: data <= 8'hFF;
            15'd733: data <= 8'hFF;
            15'd734: data <= 8'hFF;
            15'd735: data <= 8'hFF;
            15'd736: data <= 8'hFF;
            15'd737: data <= 8'hFF;
            15'd738: data <= 8'hFF;
            15'd739: data <= 8'hFF;
            15'd740: data <= 8'hFF;
            15'd741: data <= 8'hFF;
            15'd742: data <= 8'hFF;
            15'd743: data <= 8'hFF;
            15'd744: data <= 8'hFF;
            15'd745: data <= 8'h80;
            15'd746: data <= 8'h00;
            15'd747: data <= 8'h00;
            15'd748: data <= 8'h00;
            15'd749: data <= 8'h00;
            15'd750: data <= 8'h00;
            15'd751: data <= 8'h00;
            15'd752: data <= 8'h00;
            15'd753: data <= 8'h00;
            15'd754: data <= 8'h01;
            15'd755: data <= 8'hFF;
            15'd756: data <= 8'hFF;
            15'd757: data <= 8'hFF;
            15'd758: data <= 8'hFF;
            15'd759: data <= 8'hFF;
            15'd760: data <= 8'hFF;
            15'd761: data <= 8'hFF;
            15'd762: data <= 8'hFF;
            15'd763: data <= 8'hFF;
            15'd764: data <= 8'hFF;
            15'd765: data <= 8'hFF;
            15'd766: data <= 8'hFF;
            15'd767: data <= 8'hFF;
            15'd768: data <= 8'hFF;
            15'd769: data <= 8'hFF;
            15'd770: data <= 8'hFF;
            15'd771: data <= 8'hFF;
            15'd772: data <= 8'hFF;
            15'd773: data <= 8'hFF;
            15'd774: data <= 8'hFF;
            15'd775: data <= 8'h80;
            15'd776: data <= 8'h00;
            15'd777: data <= 8'h00;
            15'd778: data <= 8'h00;
            15'd779: data <= 8'h00;
            15'd780: data <= 8'h00;
            15'd781: data <= 8'h00;
            15'd782: data <= 8'h00;
            15'd783: data <= 8'h00;
            15'd784: data <= 8'h01;
            15'd785: data <= 8'hFF;
            15'd786: data <= 8'hFF;
            15'd787: data <= 8'hFF;
            15'd788: data <= 8'hFF;
            15'd789: data <= 8'hFF;
            15'd790: data <= 8'hFF;
            15'd791: data <= 8'hFF;
            15'd792: data <= 8'hFF;
            15'd793: data <= 8'hFF;
            15'd794: data <= 8'hFF;
            15'd795: data <= 8'hFF;
            15'd796: data <= 8'hFF;
            15'd797: data <= 8'hFF;
            15'd798: data <= 8'hFF;
            15'd799: data <= 8'hFF;
            15'd800: data <= 8'hFF;
            15'd801: data <= 8'hFF;
            15'd802: data <= 8'hFF;
            15'd803: data <= 8'hFF;
            15'd804: data <= 8'hFF;
            15'd805: data <= 8'h80;
            15'd806: data <= 8'h00;
            15'd807: data <= 8'h00;
            15'd808: data <= 8'h00;
            15'd809: data <= 8'h00;
            15'd810: data <= 8'h00;
            15'd811: data <= 8'h00;
            15'd812: data <= 8'h00;
            15'd813: data <= 8'h00;
            15'd814: data <= 8'h01;
            15'd815: data <= 8'hFF;
            15'd816: data <= 8'hFF;
            15'd817: data <= 8'hFF;
            15'd818: data <= 8'hFF;
            15'd819: data <= 8'hFF;
            15'd820: data <= 8'hFF;
            15'd821: data <= 8'hFF;
            15'd822: data <= 8'hFF;
            15'd823: data <= 8'hFF;
            15'd824: data <= 8'hFF;
            15'd825: data <= 8'hFF;
            15'd826: data <= 8'hFF;
            15'd827: data <= 8'hFF;
            15'd828: data <= 8'hFF;
            15'd829: data <= 8'hFF;
            15'd830: data <= 8'hFF;
            15'd831: data <= 8'hFF;
            15'd832: data <= 8'hFF;
            15'd833: data <= 8'hFF;
            15'd834: data <= 8'hFF;
            15'd835: data <= 8'h80;
            15'd836: data <= 8'h00;
            15'd837: data <= 8'h00;
            15'd838: data <= 8'h00;
            15'd839: data <= 8'h00;
            15'd840: data <= 8'h00;
            15'd841: data <= 8'h00;
            15'd842: data <= 8'h00;
            15'd843: data <= 8'h00;
            15'd844: data <= 8'h01;
            15'd845: data <= 8'hFF;
            15'd846: data <= 8'hFF;
            15'd847: data <= 8'hFF;
            15'd848: data <= 8'hFF;
            15'd849: data <= 8'hFF;
            15'd850: data <= 8'hFF;
            15'd851: data <= 8'hFF;
            15'd852: data <= 8'hFF;
            15'd853: data <= 8'hFF;
            15'd854: data <= 8'hFF;
            15'd855: data <= 8'hFF;
            15'd856: data <= 8'hFF;
            15'd857: data <= 8'hFF;
            15'd858: data <= 8'hFF;
            15'd859: data <= 8'hFF;
            15'd860: data <= 8'hFF;
            15'd861: data <= 8'hFF;
            15'd862: data <= 8'hFF;
            15'd863: data <= 8'hFF;
            15'd864: data <= 8'hFF;
            15'd865: data <= 8'h80;
            15'd866: data <= 8'h00;
            15'd867: data <= 8'h00;
            15'd868: data <= 8'h00;
            15'd869: data <= 8'h00;
            15'd870: data <= 8'h00;
            15'd871: data <= 8'h00;
            15'd872: data <= 8'h00;
            15'd873: data <= 8'h00;
            15'd874: data <= 8'h01;
            15'd875: data <= 8'hFF;
            15'd876: data <= 8'hFF;
            15'd877: data <= 8'hFF;
            15'd878: data <= 8'hFF;
            15'd879: data <= 8'hFF;
            15'd880: data <= 8'hFF;
            15'd881: data <= 8'hFF;
            15'd882: data <= 8'hFF;
            15'd883: data <= 8'hFF;
            15'd884: data <= 8'hFF;
            15'd885: data <= 8'hFF;
            15'd886: data <= 8'hFF;
            15'd887: data <= 8'hFF;
            15'd888: data <= 8'hFF;
            15'd889: data <= 8'hFF;
            15'd890: data <= 8'hFF;
            15'd891: data <= 8'hFF;
            15'd892: data <= 8'hFF;
            15'd893: data <= 8'hFF;
            15'd894: data <= 8'hFF;
            15'd895: data <= 8'h80;
            15'd896: data <= 8'h00;
            15'd897: data <= 8'h00;
            15'd898: data <= 8'h00;
            15'd899: data <= 8'h00;
            15'd900: data <= 8'h00;
            15'd901: data <= 8'h00;
            15'd902: data <= 8'h00;
            15'd903: data <= 8'h00;
            15'd904: data <= 8'h01;
            15'd905: data <= 8'hFF;
            15'd906: data <= 8'hFF;
            15'd907: data <= 8'hFF;
            15'd908: data <= 8'hFF;
            15'd909: data <= 8'hFF;
            15'd910: data <= 8'hFF;
            15'd911: data <= 8'hFF;
            15'd912: data <= 8'hFF;
            15'd913: data <= 8'hFF;
            15'd914: data <= 8'hFF;
            15'd915: data <= 8'hFF;
            15'd916: data <= 8'hFF;
            15'd917: data <= 8'hFF;
            15'd918: data <= 8'hFF;
            15'd919: data <= 8'hFF;
            15'd920: data <= 8'hFF;
            15'd921: data <= 8'hFF;
            15'd922: data <= 8'hFF;
            15'd923: data <= 8'hFF;
            15'd924: data <= 8'hFF;
            15'd925: data <= 8'h80;
            15'd926: data <= 8'h00;
            15'd927: data <= 8'h00;
            15'd928: data <= 8'h00;
            15'd929: data <= 8'h00;
            15'd930: data <= 8'h00;
            15'd931: data <= 8'h00;
            15'd932: data <= 8'h00;
            15'd933: data <= 8'h00;
            15'd934: data <= 8'h01;
            15'd935: data <= 8'hFF;
            15'd936: data <= 8'hFF;
            15'd937: data <= 8'hFF;
            15'd938: data <= 8'hFF;
            15'd939: data <= 8'hFF;
            15'd940: data <= 8'hFF;
            15'd941: data <= 8'hFF;
            15'd942: data <= 8'hFF;
            15'd943: data <= 8'hFF;
            15'd944: data <= 8'hFF;
            15'd945: data <= 8'hFF;
            15'd946: data <= 8'hFF;
            15'd947: data <= 8'hFF;
            15'd948: data <= 8'hFF;
            15'd949: data <= 8'hFF;
            15'd950: data <= 8'hFF;
            15'd951: data <= 8'hFF;
            15'd952: data <= 8'hFF;
            15'd953: data <= 8'hFF;
            15'd954: data <= 8'hFF;
            15'd955: data <= 8'h80;
            15'd956: data <= 8'h00;
            15'd957: data <= 8'h00;
            15'd958: data <= 8'h00;
            15'd959: data <= 8'h00;
            15'd960: data <= 8'h00;
            15'd961: data <= 8'h00;
            15'd962: data <= 8'h00;
            15'd963: data <= 8'h00;
            15'd964: data <= 8'h01;
            15'd965: data <= 8'hFF;
            15'd966: data <= 8'hFF;
            15'd967: data <= 8'hFF;
            15'd968: data <= 8'hFF;
            15'd969: data <= 8'hFF;
            15'd970: data <= 8'hFF;
            15'd971: data <= 8'hFF;
            15'd972: data <= 8'hFF;
            15'd973: data <= 8'hFF;
            15'd974: data <= 8'hFF;
            15'd975: data <= 8'hFF;
            15'd976: data <= 8'hFF;
            15'd977: data <= 8'hFF;
            15'd978: data <= 8'hFF;
            15'd979: data <= 8'hFF;
            15'd980: data <= 8'hFF;
            15'd981: data <= 8'hFF;
            15'd982: data <= 8'hFF;
            15'd983: data <= 8'hFF;
            15'd984: data <= 8'hFF;
            15'd985: data <= 8'h80;
            15'd986: data <= 8'h00;
            15'd987: data <= 8'h00;
            15'd988: data <= 8'h00;
            15'd989: data <= 8'h00;
            15'd990: data <= 8'h00;
            15'd991: data <= 8'h00;
            15'd992: data <= 8'h00;
            15'd993: data <= 8'h00;
            15'd994: data <= 8'h01;
            15'd995: data <= 8'hFF;
            15'd996: data <= 8'hFF;
            15'd997: data <= 8'hFF;
            15'd998: data <= 8'hFF;
            15'd999: data <= 8'hFF;
            15'd1000: data <= 8'hFF;
            15'd1001: data <= 8'hFF;
            15'd1002: data <= 8'hFF;
            15'd1003: data <= 8'hFF;
            15'd1004: data <= 8'hFF;
            15'd1005: data <= 8'hFF;
            15'd1006: data <= 8'hFF;
            15'd1007: data <= 8'hFF;
            15'd1008: data <= 8'hFF;
            15'd1009: data <= 8'hFF;
            15'd1010: data <= 8'hFF;
            15'd1011: data <= 8'hFF;
            15'd1012: data <= 8'hFF;
            15'd1013: data <= 8'hFF;
            15'd1014: data <= 8'hFF;
            15'd1015: data <= 8'h80;
            15'd1016: data <= 8'h00;
            15'd1017: data <= 8'h00;
            15'd1018: data <= 8'h00;
            15'd1019: data <= 8'h00;
            15'd1020: data <= 8'h00;
            15'd1021: data <= 8'h00;
            15'd1022: data <= 8'h00;
            15'd1023: data <= 8'h00;
            15'd1024: data <= 8'h01;
            15'd1025: data <= 8'hFF;
            15'd1026: data <= 8'hFF;
            15'd1027: data <= 8'hFF;
            15'd1028: data <= 8'hFF;
            15'd1029: data <= 8'hFF;
            15'd1030: data <= 8'hFF;
            15'd1031: data <= 8'hFF;
            15'd1032: data <= 8'hFF;
            15'd1033: data <= 8'hFF;
            15'd1034: data <= 8'hFF;
            15'd1035: data <= 8'hFF;
            15'd1036: data <= 8'hFF;
            15'd1037: data <= 8'hFF;
            15'd1038: data <= 8'hFF;
            15'd1039: data <= 8'hFF;
            15'd1040: data <= 8'hFF;
            15'd1041: data <= 8'hFF;
            15'd1042: data <= 8'hFF;
            15'd1043: data <= 8'hFF;
            15'd1044: data <= 8'hFF;
            15'd1045: data <= 8'h80;
            15'd1046: data <= 8'h00;
            15'd1047: data <= 8'h00;
            15'd1048: data <= 8'h00;
            15'd1049: data <= 8'h00;
            15'd1050: data <= 8'h00;
            15'd1051: data <= 8'h00;
            15'd1052: data <= 8'h00;
            15'd1053: data <= 8'h00;
            15'd1054: data <= 8'h01;
            15'd1055: data <= 8'hFF;
            15'd1056: data <= 8'hFF;
            15'd1057: data <= 8'hFF;
            15'd1058: data <= 8'hFF;
            15'd1059: data <= 8'hFF;
            15'd1060: data <= 8'hFF;
            15'd1061: data <= 8'hFF;
            15'd1062: data <= 8'hFF;
            15'd1063: data <= 8'hFF;
            15'd1064: data <= 8'hFF;
            15'd1065: data <= 8'hFF;
            15'd1066: data <= 8'hFF;
            15'd1067: data <= 8'hFF;
            15'd1068: data <= 8'hFF;
            15'd1069: data <= 8'hFF;
            15'd1070: data <= 8'hFF;
            15'd1071: data <= 8'hFF;
            15'd1072: data <= 8'hFF;
            15'd1073: data <= 8'hFF;
            15'd1074: data <= 8'hFF;
            15'd1075: data <= 8'h80;
            15'd1076: data <= 8'h00;
            15'd1077: data <= 8'h00;
            15'd1078: data <= 8'h00;
            15'd1079: data <= 8'h00;
            15'd1080: data <= 8'h00;
            15'd1081: data <= 8'h00;
            15'd1082: data <= 8'h00;
            15'd1083: data <= 8'h00;
            15'd1084: data <= 8'h01;
            15'd1085: data <= 8'hFF;
            15'd1086: data <= 8'hFF;
            15'd1087: data <= 8'hFF;
            15'd1088: data <= 8'hFF;
            15'd1089: data <= 8'hFF;
            15'd1090: data <= 8'hFF;
            15'd1091: data <= 8'hFF;
            15'd1092: data <= 8'hFF;
            15'd1093: data <= 8'hFF;
            15'd1094: data <= 8'hFF;
            15'd1095: data <= 8'hFF;
            15'd1096: data <= 8'hFF;
            15'd1097: data <= 8'hFF;
            15'd1098: data <= 8'hFF;
            15'd1099: data <= 8'hFF;
            15'd1100: data <= 8'hFF;
            15'd1101: data <= 8'hFF;
            15'd1102: data <= 8'hFF;
            15'd1103: data <= 8'hFF;
            15'd1104: data <= 8'hFF;
            15'd1105: data <= 8'h80;
            15'd1106: data <= 8'h00;
            15'd1107: data <= 8'h00;
            15'd1108: data <= 8'h00;
            15'd1109: data <= 8'h00;
            15'd1110: data <= 8'h00;
            15'd1111: data <= 8'h00;
            15'd1112: data <= 8'h00;
            15'd1113: data <= 8'h00;
            15'd1114: data <= 8'h01;
            15'd1115: data <= 8'hFF;
            15'd1116: data <= 8'hFF;
            15'd1117: data <= 8'hFF;
            15'd1118: data <= 8'hFF;
            15'd1119: data <= 8'hFF;
            15'd1120: data <= 8'hFF;
            15'd1121: data <= 8'hFF;
            15'd1122: data <= 8'hFF;
            15'd1123: data <= 8'hFF;
            15'd1124: data <= 8'hFF;
            15'd1125: data <= 8'hFF;
            15'd1126: data <= 8'hFF;
            15'd1127: data <= 8'hFF;
            15'd1128: data <= 8'hFF;
            15'd1129: data <= 8'hFF;
            15'd1130: data <= 8'hFF;
            15'd1131: data <= 8'hFF;
            15'd1132: data <= 8'hFF;
            15'd1133: data <= 8'hFF;
            15'd1134: data <= 8'hFF;
            15'd1135: data <= 8'h80;
            15'd1136: data <= 8'h00;
            15'd1137: data <= 8'h00;
            15'd1138: data <= 8'h00;
            15'd1139: data <= 8'h00;
            15'd1140: data <= 8'h00;
            15'd1141: data <= 8'h00;
            15'd1142: data <= 8'h00;
            15'd1143: data <= 8'h00;
            15'd1144: data <= 8'h01;
            15'd1145: data <= 8'hFF;
            15'd1146: data <= 8'hFF;
            15'd1147: data <= 8'hFF;
            15'd1148: data <= 8'hFF;
            15'd1149: data <= 8'hFF;
            15'd1150: data <= 8'hFF;
            15'd1151: data <= 8'hFF;
            15'd1152: data <= 8'hFF;
            15'd1153: data <= 8'hFF;
            15'd1154: data <= 8'hFF;
            15'd1155: data <= 8'hFF;
            15'd1156: data <= 8'hFF;
            15'd1157: data <= 8'hFF;
            15'd1158: data <= 8'hFF;
            15'd1159: data <= 8'hFF;
            15'd1160: data <= 8'hFF;
            15'd1161: data <= 8'hFF;
            15'd1162: data <= 8'hFF;
            15'd1163: data <= 8'hFF;
            15'd1164: data <= 8'hFF;
            15'd1165: data <= 8'h80;
            15'd1166: data <= 8'h00;
            15'd1167: data <= 8'h00;
            15'd1168: data <= 8'h00;
            15'd1169: data <= 8'h00;
            15'd1170: data <= 8'h00;
            15'd1171: data <= 8'h00;
            15'd1172: data <= 8'h00;
            15'd1173: data <= 8'h00;
            15'd1174: data <= 8'h01;
            15'd1175: data <= 8'hFF;
            15'd1176: data <= 8'hFF;
            15'd1177: data <= 8'hFF;
            15'd1178: data <= 8'hFF;
            15'd1179: data <= 8'hFF;
            15'd1180: data <= 8'hFF;
            15'd1181: data <= 8'hFF;
            15'd1182: data <= 8'hFF;
            15'd1183: data <= 8'hFF;
            15'd1184: data <= 8'hFF;
            15'd1185: data <= 8'hFF;
            15'd1186: data <= 8'hFF;
            15'd1187: data <= 8'hFF;
            15'd1188: data <= 8'hFF;
            15'd1189: data <= 8'hFF;
            15'd1190: data <= 8'hFF;
            15'd1191: data <= 8'hFF;
            15'd1192: data <= 8'hFF;
            15'd1193: data <= 8'hFF;
            15'd1194: data <= 8'hFF;
            15'd1195: data <= 8'h80;
            15'd1196: data <= 8'h00;
            15'd1197: data <= 8'h00;
            15'd1198: data <= 8'h00;
            15'd1199: data <= 8'h00;
            15'd1200: data <= 8'h00;
            15'd1201: data <= 8'h00;
            15'd1202: data <= 8'h00;
            15'd1203: data <= 8'h00;
            15'd1204: data <= 8'h01;
            15'd1205: data <= 8'hFF;
            15'd1206: data <= 8'hFF;
            15'd1207: data <= 8'hFF;
            15'd1208: data <= 8'hFF;
            15'd1209: data <= 8'hFF;
            15'd1210: data <= 8'hFF;
            15'd1211: data <= 8'hFF;
            15'd1212: data <= 8'hFF;
            15'd1213: data <= 8'hFF;
            15'd1214: data <= 8'hFF;
            15'd1215: data <= 8'hFF;
            15'd1216: data <= 8'hFF;
            15'd1217: data <= 8'hFF;
            15'd1218: data <= 8'hFF;
            15'd1219: data <= 8'hFF;
            15'd1220: data <= 8'hFF;
            15'd1221: data <= 8'hFF;
            15'd1222: data <= 8'hFF;
            15'd1223: data <= 8'hFF;
            15'd1224: data <= 8'hFF;
            15'd1225: data <= 8'h80;
            15'd1226: data <= 8'h00;
            15'd1227: data <= 8'h00;
            15'd1228: data <= 8'h00;
            15'd1229: data <= 8'h00;
            15'd1230: data <= 8'h00;
            15'd1231: data <= 8'h00;
            15'd1232: data <= 8'h00;
            15'd1233: data <= 8'h00;
            15'd1234: data <= 8'h01;
            15'd1235: data <= 8'hFF;
            15'd1236: data <= 8'hFF;
            15'd1237: data <= 8'hFF;
            15'd1238: data <= 8'hFF;
            15'd1239: data <= 8'hFF;
            15'd1240: data <= 8'hFF;
            15'd1241: data <= 8'hFF;
            15'd1242: data <= 8'hFF;
            15'd1243: data <= 8'hFF;
            15'd1244: data <= 8'hFF;
            15'd1245: data <= 8'hFF;
            15'd1246: data <= 8'hFF;
            15'd1247: data <= 8'hFF;
            15'd1248: data <= 8'hFF;
            15'd1249: data <= 8'hFF;
            15'd1250: data <= 8'hFF;
            15'd1251: data <= 8'hFF;
            15'd1252: data <= 8'hFF;
            15'd1253: data <= 8'hFF;
            15'd1254: data <= 8'hFF;
            15'd1255: data <= 8'h80;
            15'd1256: data <= 8'h00;
            15'd1257: data <= 8'h00;
            15'd1258: data <= 8'h00;
            15'd1259: data <= 8'h00;
            15'd1260: data <= 8'h00;
            15'd1261: data <= 8'h00;
            15'd1262: data <= 8'h00;
            15'd1263: data <= 8'h00;
            15'd1264: data <= 8'h01;
            15'd1265: data <= 8'hFF;
            15'd1266: data <= 8'hFF;
            15'd1267: data <= 8'hFF;
            15'd1268: data <= 8'hFF;
            15'd1269: data <= 8'hFF;
            15'd1270: data <= 8'hFF;
            15'd1271: data <= 8'hFF;
            15'd1272: data <= 8'hFF;
            15'd1273: data <= 8'hFF;
            15'd1274: data <= 8'hFF;
            15'd1275: data <= 8'hFF;
            15'd1276: data <= 8'hFF;
            15'd1277: data <= 8'hFF;
            15'd1278: data <= 8'hFF;
            15'd1279: data <= 8'hFF;
            15'd1280: data <= 8'hFF;
            15'd1281: data <= 8'hFF;
            15'd1282: data <= 8'hFF;
            15'd1283: data <= 8'hFF;
            15'd1284: data <= 8'hFF;
            15'd1285: data <= 8'h80;
            15'd1286: data <= 8'h00;
            15'd1287: data <= 8'h00;
            15'd1288: data <= 8'h00;
            15'd1289: data <= 8'h00;
            15'd1290: data <= 8'h00;
            15'd1291: data <= 8'h00;
            15'd1292: data <= 8'h00;
            15'd1293: data <= 8'h00;
            15'd1294: data <= 8'h01;
            15'd1295: data <= 8'hFF;
            15'd1296: data <= 8'hFF;
            15'd1297: data <= 8'hFF;
            15'd1298: data <= 8'hFF;
            15'd1299: data <= 8'hFF;
            15'd1300: data <= 8'hFF;
            15'd1301: data <= 8'hFF;
            15'd1302: data <= 8'hFF;
            15'd1303: data <= 8'hFF;
            15'd1304: data <= 8'hFF;
            15'd1305: data <= 8'hFF;
            15'd1306: data <= 8'hFF;
            15'd1307: data <= 8'hFF;
            15'd1308: data <= 8'hFF;
            15'd1309: data <= 8'hFF;
            15'd1310: data <= 8'hFF;
            15'd1311: data <= 8'hFF;
            15'd1312: data <= 8'hFF;
            15'd1313: data <= 8'hFF;
            15'd1314: data <= 8'hFF;
            15'd1315: data <= 8'h80;
            15'd1316: data <= 8'h00;
            15'd1317: data <= 8'h00;
            15'd1318: data <= 8'h00;
            15'd1319: data <= 8'h00;
            15'd1320: data <= 8'h00;
            15'd1321: data <= 8'h00;
            15'd1322: data <= 8'h00;
            15'd1323: data <= 8'h00;
            15'd1324: data <= 8'h01;
            15'd1325: data <= 8'hFF;
            15'd1326: data <= 8'hFF;
            15'd1327: data <= 8'hFF;
            15'd1328: data <= 8'hFF;
            15'd1329: data <= 8'hFF;
            15'd1330: data <= 8'hFF;
            15'd1331: data <= 8'hFF;
            15'd1332: data <= 8'hFF;
            15'd1333: data <= 8'hFF;
            15'd1334: data <= 8'hFF;
            15'd1335: data <= 8'hFF;
            15'd1336: data <= 8'hFF;
            15'd1337: data <= 8'hFF;
            15'd1338: data <= 8'hFF;
            15'd1339: data <= 8'hFF;
            15'd1340: data <= 8'hFF;
            15'd1341: data <= 8'hFF;
            15'd1342: data <= 8'hFF;
            15'd1343: data <= 8'hFF;
            15'd1344: data <= 8'hFF;
            15'd1345: data <= 8'h80;
            15'd1346: data <= 8'h00;
            15'd1347: data <= 8'h00;
            15'd1348: data <= 8'h00;
            15'd1349: data <= 8'h00;
            15'd1350: data <= 8'h00;
            15'd1351: data <= 8'h00;
            15'd1352: data <= 8'h00;
            15'd1353: data <= 8'h00;
            15'd1354: data <= 8'h01;
            15'd1355: data <= 8'hFF;
            15'd1356: data <= 8'hFF;
            15'd1357: data <= 8'hFF;
            15'd1358: data <= 8'hFF;
            15'd1359: data <= 8'hFF;
            15'd1360: data <= 8'hFF;
            15'd1361: data <= 8'hFF;
            15'd1362: data <= 8'hFF;
            15'd1363: data <= 8'hFF;
            15'd1364: data <= 8'hFF;
            15'd1365: data <= 8'hFF;
            15'd1366: data <= 8'hFF;
            15'd1367: data <= 8'hFF;
            15'd1368: data <= 8'hFF;
            15'd1369: data <= 8'hFF;
            15'd1370: data <= 8'hFF;
            15'd1371: data <= 8'hFF;
            15'd1372: data <= 8'hFF;
            15'd1373: data <= 8'hFF;
            15'd1374: data <= 8'hFF;
            15'd1375: data <= 8'h80;
            15'd1376: data <= 8'h00;
            15'd1377: data <= 8'h00;
            15'd1378: data <= 8'h00;
            15'd1379: data <= 8'h00;
            15'd1380: data <= 8'h00;
            15'd1381: data <= 8'h00;
            15'd1382: data <= 8'h00;
            15'd1383: data <= 8'h00;
            15'd1384: data <= 8'h01;
            15'd1385: data <= 8'hFF;
            15'd1386: data <= 8'hFF;
            15'd1387: data <= 8'hFF;
            15'd1388: data <= 8'hFF;
            15'd1389: data <= 8'hFF;
            15'd1390: data <= 8'hFF;
            15'd1391: data <= 8'hFF;
            15'd1392: data <= 8'hFF;
            15'd1393: data <= 8'hFF;
            15'd1394: data <= 8'hFF;
            15'd1395: data <= 8'hFF;
            15'd1396: data <= 8'hFF;
            15'd1397: data <= 8'hF7;
            15'd1398: data <= 8'hFF;
            15'd1399: data <= 8'hFF;
            15'd1400: data <= 8'hFF;
            15'd1401: data <= 8'hFF;
            15'd1402: data <= 8'hFF;
            15'd1403: data <= 8'hFF;
            15'd1404: data <= 8'hFF;
            15'd1405: data <= 8'h80;
            15'd1406: data <= 8'h00;
            15'd1407: data <= 8'h00;
            15'd1408: data <= 8'h00;
            15'd1409: data <= 8'h00;
            15'd1410: data <= 8'h00;
            15'd1411: data <= 8'h00;
            15'd1412: data <= 8'h00;
            15'd1413: data <= 8'h00;
            15'd1414: data <= 8'h01;
            15'd1415: data <= 8'hFF;
            15'd1416: data <= 8'hFF;
            15'd1417: data <= 8'hFF;
            15'd1418: data <= 8'hFF;
            15'd1419: data <= 8'hFF;
            15'd1420: data <= 8'hFF;
            15'd1421: data <= 8'hFF;
            15'd1422: data <= 8'h83;
            15'd1423: data <= 8'hFF;
            15'd1424: data <= 8'hFF;
            15'd1425: data <= 8'hFF;
            15'd1426: data <= 8'hFF;
            15'd1427: data <= 8'h03;
            15'd1428: data <= 8'hFF;
            15'd1429: data <= 8'hFF;
            15'd1430: data <= 8'hFF;
            15'd1431: data <= 8'hFF;
            15'd1432: data <= 8'hFF;
            15'd1433: data <= 8'hFF;
            15'd1434: data <= 8'hFF;
            15'd1435: data <= 8'h80;
            15'd1436: data <= 8'h00;
            15'd1437: data <= 8'h00;
            15'd1438: data <= 8'h00;
            15'd1439: data <= 8'h00;
            15'd1440: data <= 8'h00;
            15'd1441: data <= 8'h00;
            15'd1442: data <= 8'h00;
            15'd1443: data <= 8'h00;
            15'd1444: data <= 8'h01;
            15'd1445: data <= 8'hFF;
            15'd1446: data <= 8'hFF;
            15'd1447: data <= 8'hFF;
            15'd1448: data <= 8'hFF;
            15'd1449: data <= 8'hFF;
            15'd1450: data <= 8'hFF;
            15'd1451: data <= 8'hFF;
            15'd1452: data <= 8'h80;
            15'd1453: data <= 8'h7F;
            15'd1454: data <= 8'hFF;
            15'd1455: data <= 8'hFF;
            15'd1456: data <= 8'hFC;
            15'd1457: data <= 8'h03;
            15'd1458: data <= 8'hFF;
            15'd1459: data <= 8'hFF;
            15'd1460: data <= 8'hFF;
            15'd1461: data <= 8'hFF;
            15'd1462: data <= 8'hFF;
            15'd1463: data <= 8'hFF;
            15'd1464: data <= 8'hFF;
            15'd1465: data <= 8'h80;
            15'd1466: data <= 8'h00;
            15'd1467: data <= 8'h00;
            15'd1468: data <= 8'h00;
            15'd1469: data <= 8'h00;
            15'd1470: data <= 8'h00;
            15'd1471: data <= 8'h00;
            15'd1472: data <= 8'h00;
            15'd1473: data <= 8'h00;
            15'd1474: data <= 8'h01;
            15'd1475: data <= 8'hFF;
            15'd1476: data <= 8'hFF;
            15'd1477: data <= 8'hFF;
            15'd1478: data <= 8'hFF;
            15'd1479: data <= 8'hFF;
            15'd1480: data <= 8'hFF;
            15'd1481: data <= 8'hFF;
            15'd1482: data <= 8'h00;
            15'd1483: data <= 8'h07;
            15'd1484: data <= 8'hFF;
            15'd1485: data <= 8'hFF;
            15'd1486: data <= 8'hF8;
            15'd1487: data <= 8'h03;
            15'd1488: data <= 8'hFF;
            15'd1489: data <= 8'hFF;
            15'd1490: data <= 8'hFF;
            15'd1491: data <= 8'hFF;
            15'd1492: data <= 8'hFF;
            15'd1493: data <= 8'hFF;
            15'd1494: data <= 8'hFF;
            15'd1495: data <= 8'h80;
            15'd1496: data <= 8'h00;
            15'd1497: data <= 8'h00;
            15'd1498: data <= 8'h00;
            15'd1499: data <= 8'h00;
            15'd1500: data <= 8'h00;
            15'd1501: data <= 8'h00;
            15'd1502: data <= 8'h00;
            15'd1503: data <= 8'h00;
            15'd1504: data <= 8'h01;
            15'd1505: data <= 8'hFF;
            15'd1506: data <= 8'hFF;
            15'd1507: data <= 8'hFF;
            15'd1508: data <= 8'hFF;
            15'd1509: data <= 8'hFF;
            15'd1510: data <= 8'hFF;
            15'd1511: data <= 8'hFF;
            15'd1512: data <= 8'h80;
            15'd1513: data <= 8'h01;
            15'd1514: data <= 8'hFF;
            15'd1515: data <= 8'hFF;
            15'd1516: data <= 8'hE0;
            15'd1517: data <= 8'h07;
            15'd1518: data <= 8'hFF;
            15'd1519: data <= 8'hFF;
            15'd1520: data <= 8'hFF;
            15'd1521: data <= 8'hFF;
            15'd1522: data <= 8'hFF;
            15'd1523: data <= 8'hFF;
            15'd1524: data <= 8'hFF;
            15'd1525: data <= 8'h80;
            15'd1526: data <= 8'h00;
            15'd1527: data <= 8'h00;
            15'd1528: data <= 8'h00;
            15'd1529: data <= 8'h00;
            15'd1530: data <= 8'h00;
            15'd1531: data <= 8'h00;
            15'd1532: data <= 8'h00;
            15'd1533: data <= 8'h00;
            15'd1534: data <= 8'h01;
            15'd1535: data <= 8'hFF;
            15'd1536: data <= 8'hFF;
            15'd1537: data <= 8'hFF;
            15'd1538: data <= 8'hFF;
            15'd1539: data <= 8'hFF;
            15'd1540: data <= 8'hFF;
            15'd1541: data <= 8'hFF;
            15'd1542: data <= 8'hE0;
            15'd1543: data <= 8'h00;
            15'd1544: data <= 8'hFF;
            15'd1545: data <= 8'hFF;
            15'd1546: data <= 8'hC0;
            15'd1547: data <= 8'h1F;
            15'd1548: data <= 8'hFF;
            15'd1549: data <= 8'hFF;
            15'd1550: data <= 8'hFF;
            15'd1551: data <= 8'hFF;
            15'd1552: data <= 8'hFF;
            15'd1553: data <= 8'hFF;
            15'd1554: data <= 8'hFF;
            15'd1555: data <= 8'h80;
            15'd1556: data <= 8'h00;
            15'd1557: data <= 8'h00;
            15'd1558: data <= 8'h00;
            15'd1559: data <= 8'h00;
            15'd1560: data <= 8'h00;
            15'd1561: data <= 8'h00;
            15'd1562: data <= 8'h00;
            15'd1563: data <= 8'h00;
            15'd1564: data <= 8'h01;
            15'd1565: data <= 8'hFF;
            15'd1566: data <= 8'hFF;
            15'd1567: data <= 8'hFF;
            15'd1568: data <= 8'hFF;
            15'd1569: data <= 8'hFF;
            15'd1570: data <= 8'hFF;
            15'd1571: data <= 8'hFF;
            15'd1572: data <= 8'hFC;
            15'd1573: data <= 8'h00;
            15'd1574: data <= 8'h7F;
            15'd1575: data <= 8'hFF;
            15'd1576: data <= 8'h00;
            15'd1577: data <= 8'h7F;
            15'd1578: data <= 8'hFF;
            15'd1579: data <= 8'hFF;
            15'd1580: data <= 8'hFF;
            15'd1581: data <= 8'hFF;
            15'd1582: data <= 8'hFF;
            15'd1583: data <= 8'hFF;
            15'd1584: data <= 8'hFF;
            15'd1585: data <= 8'h80;
            15'd1586: data <= 8'h00;
            15'd1587: data <= 8'h00;
            15'd1588: data <= 8'h00;
            15'd1589: data <= 8'h00;
            15'd1590: data <= 8'h00;
            15'd1591: data <= 8'h00;
            15'd1592: data <= 8'h00;
            15'd1593: data <= 8'h00;
            15'd1594: data <= 8'h01;
            15'd1595: data <= 8'hFF;
            15'd1596: data <= 8'hFF;
            15'd1597: data <= 8'hFF;
            15'd1598: data <= 8'hFF;
            15'd1599: data <= 8'hFF;
            15'd1600: data <= 8'hFF;
            15'd1601: data <= 8'hFF;
            15'd1602: data <= 8'hFF;
            15'd1603: data <= 8'h00;
            15'd1604: data <= 8'hFF;
            15'd1605: data <= 8'hFF;
            15'd1606: data <= 8'h01;
            15'd1607: data <= 8'hFF;
            15'd1608: data <= 8'hFF;
            15'd1609: data <= 8'hFF;
            15'd1610: data <= 8'hFF;
            15'd1611: data <= 8'hFF;
            15'd1612: data <= 8'hFF;
            15'd1613: data <= 8'hFF;
            15'd1614: data <= 8'hFF;
            15'd1615: data <= 8'h80;
            15'd1616: data <= 8'h00;
            15'd1617: data <= 8'h00;
            15'd1618: data <= 8'h00;
            15'd1619: data <= 8'h00;
            15'd1620: data <= 8'h00;
            15'd1621: data <= 8'h00;
            15'd1622: data <= 8'h00;
            15'd1623: data <= 8'h00;
            15'd1624: data <= 8'h01;
            15'd1625: data <= 8'hFF;
            15'd1626: data <= 8'hFF;
            15'd1627: data <= 8'hFF;
            15'd1628: data <= 8'hFF;
            15'd1629: data <= 8'hFF;
            15'd1630: data <= 8'hFF;
            15'd1631: data <= 8'hFF;
            15'd1632: data <= 8'hFF;
            15'd1633: data <= 8'hF1;
            15'd1634: data <= 8'hFF;
            15'd1635: data <= 8'hFE;
            15'd1636: data <= 8'h07;
            15'd1637: data <= 8'hFF;
            15'd1638: data <= 8'hFF;
            15'd1639: data <= 8'hFF;
            15'd1640: data <= 8'hFF;
            15'd1641: data <= 8'hFF;
            15'd1642: data <= 8'hFF;
            15'd1643: data <= 8'hFF;
            15'd1644: data <= 8'hFF;
            15'd1645: data <= 8'h80;
            15'd1646: data <= 8'h00;
            15'd1647: data <= 8'h00;
            15'd1648: data <= 8'h00;
            15'd1649: data <= 8'h00;
            15'd1650: data <= 8'h00;
            15'd1651: data <= 8'h00;
            15'd1652: data <= 8'h00;
            15'd1653: data <= 8'h00;
            15'd1654: data <= 8'h01;
            15'd1655: data <= 8'hFF;
            15'd1656: data <= 8'hFF;
            15'd1657: data <= 8'hFF;
            15'd1658: data <= 8'hFF;
            15'd1659: data <= 8'hFF;
            15'd1660: data <= 8'hFF;
            15'd1661: data <= 8'hFF;
            15'd1662: data <= 8'hFF;
            15'd1663: data <= 8'hFF;
            15'd1664: data <= 8'hFF;
            15'd1665: data <= 8'hFF;
            15'd1666: data <= 8'h1F;
            15'd1667: data <= 8'hFF;
            15'd1668: data <= 8'hFF;
            15'd1669: data <= 8'hFF;
            15'd1670: data <= 8'hFF;
            15'd1671: data <= 8'hFF;
            15'd1672: data <= 8'hFF;
            15'd1673: data <= 8'hFF;
            15'd1674: data <= 8'hFF;
            15'd1675: data <= 8'h80;
            15'd1676: data <= 8'h00;
            15'd1677: data <= 8'h00;
            15'd1678: data <= 8'h00;
            15'd1679: data <= 8'h00;
            15'd1680: data <= 8'h00;
            15'd1681: data <= 8'h00;
            15'd1682: data <= 8'h00;
            15'd1683: data <= 8'h00;
            15'd1684: data <= 8'h01;
            15'd1685: data <= 8'hFF;
            15'd1686: data <= 8'hFF;
            15'd1687: data <= 8'hFF;
            15'd1688: data <= 8'hFF;
            15'd1689: data <= 8'hFF;
            15'd1690: data <= 8'hFF;
            15'd1691: data <= 8'hFF;
            15'd1692: data <= 8'hFF;
            15'd1693: data <= 8'hFF;
            15'd1694: data <= 8'hFF;
            15'd1695: data <= 8'hFF;
            15'd1696: data <= 8'hFF;
            15'd1697: data <= 8'hFF;
            15'd1698: data <= 8'hFF;
            15'd1699: data <= 8'hFF;
            15'd1700: data <= 8'hFF;
            15'd1701: data <= 8'hFF;
            15'd1702: data <= 8'hFF;
            15'd1703: data <= 8'hFF;
            15'd1704: data <= 8'hFF;
            15'd1705: data <= 8'h80;
            15'd1706: data <= 8'h00;
            15'd1707: data <= 8'h00;
            15'd1708: data <= 8'h00;
            15'd1709: data <= 8'h00;
            15'd1710: data <= 8'h00;
            15'd1711: data <= 8'h00;
            15'd1712: data <= 8'h00;
            15'd1713: data <= 8'h00;
            15'd1714: data <= 8'h01;
            15'd1715: data <= 8'hFF;
            15'd1716: data <= 8'hFF;
            15'd1717: data <= 8'hFF;
            15'd1718: data <= 8'hFF;
            15'd1719: data <= 8'hFF;
            15'd1720: data <= 8'hFF;
            15'd1721: data <= 8'hFF;
            15'd1722: data <= 8'hFF;
            15'd1723: data <= 8'hFF;
            15'd1724: data <= 8'hFF;
            15'd1725: data <= 8'hFF;
            15'd1726: data <= 8'hFF;
            15'd1727: data <= 8'hFF;
            15'd1728: data <= 8'hFF;
            15'd1729: data <= 8'hFF;
            15'd1730: data <= 8'hFF;
            15'd1731: data <= 8'hFF;
            15'd1732: data <= 8'hFF;
            15'd1733: data <= 8'hFF;
            15'd1734: data <= 8'hFF;
            15'd1735: data <= 8'h80;
            15'd1736: data <= 8'h00;
            15'd1737: data <= 8'h00;
            15'd1738: data <= 8'h00;
            15'd1739: data <= 8'h00;
            15'd1740: data <= 8'h00;
            15'd1741: data <= 8'h00;
            15'd1742: data <= 8'h00;
            15'd1743: data <= 8'h00;
            15'd1744: data <= 8'h01;
            15'd1745: data <= 8'hFF;
            15'd1746: data <= 8'hFF;
            15'd1747: data <= 8'hFF;
            15'd1748: data <= 8'hFF;
            15'd1749: data <= 8'hFF;
            15'd1750: data <= 8'hFF;
            15'd1751: data <= 8'hFF;
            15'd1752: data <= 8'hFF;
            15'd1753: data <= 8'hDF;
            15'd1754: data <= 8'hFF;
            15'd1755: data <= 8'hFF;
            15'd1756: data <= 8'hFF;
            15'd1757: data <= 8'hFF;
            15'd1758: data <= 8'hFF;
            15'd1759: data <= 8'hFF;
            15'd1760: data <= 8'hFF;
            15'd1761: data <= 8'hFF;
            15'd1762: data <= 8'hFF;
            15'd1763: data <= 8'hFF;
            15'd1764: data <= 8'hFF;
            15'd1765: data <= 8'h80;
            15'd1766: data <= 8'h00;
            15'd1767: data <= 8'h00;
            15'd1768: data <= 8'h00;
            15'd1769: data <= 8'h00;
            15'd1770: data <= 8'h00;
            15'd1771: data <= 8'h00;
            15'd1772: data <= 8'h00;
            15'd1773: data <= 8'h00;
            15'd1774: data <= 8'h01;
            15'd1775: data <= 8'hFF;
            15'd1776: data <= 8'hFF;
            15'd1777: data <= 8'hFF;
            15'd1778: data <= 8'hFF;
            15'd1779: data <= 8'hFF;
            15'd1780: data <= 8'hFF;
            15'd1781: data <= 8'hFF;
            15'd1782: data <= 8'hFF;
            15'd1783: data <= 8'h07;
            15'd1784: data <= 8'hFF;
            15'd1785: data <= 8'hFF;
            15'd1786: data <= 8'hF0;
            15'd1787: data <= 8'h7F;
            15'd1788: data <= 8'hFF;
            15'd1789: data <= 8'hFF;
            15'd1790: data <= 8'hFF;
            15'd1791: data <= 8'hFF;
            15'd1792: data <= 8'hFF;
            15'd1793: data <= 8'hFF;
            15'd1794: data <= 8'hFF;
            15'd1795: data <= 8'h80;
            15'd1796: data <= 8'h00;
            15'd1797: data <= 8'h00;
            15'd1798: data <= 8'h00;
            15'd1799: data <= 8'h00;
            15'd1800: data <= 8'h00;
            15'd1801: data <= 8'h00;
            15'd1802: data <= 8'h00;
            15'd1803: data <= 8'h00;
            15'd1804: data <= 8'h01;
            15'd1805: data <= 8'hFF;
            15'd1806: data <= 8'hFF;
            15'd1807: data <= 8'hFF;
            15'd1808: data <= 8'hFF;
            15'd1809: data <= 8'hFF;
            15'd1810: data <= 8'hFF;
            15'd1811: data <= 8'hFF;
            15'd1812: data <= 8'hFE;
            15'd1813: data <= 8'h07;
            15'd1814: data <= 8'hFF;
            15'd1815: data <= 8'hFF;
            15'd1816: data <= 8'hE0;
            15'd1817: data <= 8'h7F;
            15'd1818: data <= 8'hFF;
            15'd1819: data <= 8'hFF;
            15'd1820: data <= 8'hFF;
            15'd1821: data <= 8'hFF;
            15'd1822: data <= 8'hFF;
            15'd1823: data <= 8'hFF;
            15'd1824: data <= 8'hFF;
            15'd1825: data <= 8'h80;
            15'd1826: data <= 8'h00;
            15'd1827: data <= 8'h00;
            15'd1828: data <= 8'h00;
            15'd1829: data <= 8'h00;
            15'd1830: data <= 8'h00;
            15'd1831: data <= 8'h00;
            15'd1832: data <= 8'h00;
            15'd1833: data <= 8'h00;
            15'd1834: data <= 8'h01;
            15'd1835: data <= 8'hFF;
            15'd1836: data <= 8'hFF;
            15'd1837: data <= 8'hFF;
            15'd1838: data <= 8'hFF;
            15'd1839: data <= 8'hFF;
            15'd1840: data <= 8'hFF;
            15'd1841: data <= 8'hFF;
            15'd1842: data <= 8'hFC;
            15'd1843: data <= 8'h03;
            15'd1844: data <= 8'hFF;
            15'd1845: data <= 8'hFF;
            15'd1846: data <= 8'hC0;
            15'd1847: data <= 8'h3F;
            15'd1848: data <= 8'hFF;
            15'd1849: data <= 8'hFF;
            15'd1850: data <= 8'hFF;
            15'd1851: data <= 8'hFF;
            15'd1852: data <= 8'hFF;
            15'd1853: data <= 8'hFF;
            15'd1854: data <= 8'hFF;
            15'd1855: data <= 8'h80;
            15'd1856: data <= 8'h00;
            15'd1857: data <= 8'h00;
            15'd1858: data <= 8'h00;
            15'd1859: data <= 8'h00;
            15'd1860: data <= 8'h00;
            15'd1861: data <= 8'h00;
            15'd1862: data <= 8'h00;
            15'd1863: data <= 8'h00;
            15'd1864: data <= 8'h01;
            15'd1865: data <= 8'hFF;
            15'd1866: data <= 8'hFF;
            15'd1867: data <= 8'hFF;
            15'd1868: data <= 8'hFF;
            15'd1869: data <= 8'hFF;
            15'd1870: data <= 8'hFF;
            15'd1871: data <= 8'hFF;
            15'd1872: data <= 8'hFC;
            15'd1873: data <= 8'h03;
            15'd1874: data <= 8'hFF;
            15'd1875: data <= 8'hFF;
            15'd1876: data <= 8'hC0;
            15'd1877: data <= 8'h3F;
            15'd1878: data <= 8'hFF;
            15'd1879: data <= 8'hFF;
            15'd1880: data <= 8'hFF;
            15'd1881: data <= 8'hFF;
            15'd1882: data <= 8'hFF;
            15'd1883: data <= 8'hFF;
            15'd1884: data <= 8'hFF;
            15'd1885: data <= 8'h80;
            15'd1886: data <= 8'h00;
            15'd1887: data <= 8'h00;
            15'd1888: data <= 8'h00;
            15'd1889: data <= 8'h00;
            15'd1890: data <= 8'h00;
            15'd1891: data <= 8'h00;
            15'd1892: data <= 8'h00;
            15'd1893: data <= 8'h00;
            15'd1894: data <= 8'h01;
            15'd1895: data <= 8'hFF;
            15'd1896: data <= 8'hFF;
            15'd1897: data <= 8'hFF;
            15'd1898: data <= 8'hFF;
            15'd1899: data <= 8'hFF;
            15'd1900: data <= 8'hFF;
            15'd1901: data <= 8'hFF;
            15'd1902: data <= 8'hFC;
            15'd1903: data <= 8'h03;
            15'd1904: data <= 8'hFF;
            15'd1905: data <= 8'hFF;
            15'd1906: data <= 8'hC0;
            15'd1907: data <= 8'h3F;
            15'd1908: data <= 8'hFF;
            15'd1909: data <= 8'hFF;
            15'd1910: data <= 8'hFF;
            15'd1911: data <= 8'hFF;
            15'd1912: data <= 8'hFF;
            15'd1913: data <= 8'hFF;
            15'd1914: data <= 8'hFF;
            15'd1915: data <= 8'h80;
            15'd1916: data <= 8'h00;
            15'd1917: data <= 8'h00;
            15'd1918: data <= 8'h00;
            15'd1919: data <= 8'h00;
            15'd1920: data <= 8'h00;
            15'd1921: data <= 8'h00;
            15'd1922: data <= 8'h00;
            15'd1923: data <= 8'h00;
            15'd1924: data <= 8'h01;
            15'd1925: data <= 8'hFF;
            15'd1926: data <= 8'hFF;
            15'd1927: data <= 8'hFF;
            15'd1928: data <= 8'hFF;
            15'd1929: data <= 8'hFF;
            15'd1930: data <= 8'hFF;
            15'd1931: data <= 8'hFF;
            15'd1932: data <= 8'hFC;
            15'd1933: data <= 8'h03;
            15'd1934: data <= 8'hFF;
            15'd1935: data <= 8'hFF;
            15'd1936: data <= 8'hC0;
            15'd1937: data <= 8'h7F;
            15'd1938: data <= 8'hFF;
            15'd1939: data <= 8'hFF;
            15'd1940: data <= 8'hFF;
            15'd1941: data <= 8'hFF;
            15'd1942: data <= 8'hFF;
            15'd1943: data <= 8'hFF;
            15'd1944: data <= 8'hFF;
            15'd1945: data <= 8'h80;
            15'd1946: data <= 8'h00;
            15'd1947: data <= 8'h00;
            15'd1948: data <= 8'h00;
            15'd1949: data <= 8'h00;
            15'd1950: data <= 8'h00;
            15'd1951: data <= 8'h00;
            15'd1952: data <= 8'h00;
            15'd1953: data <= 8'h00;
            15'd1954: data <= 8'h01;
            15'd1955: data <= 8'hFF;
            15'd1956: data <= 8'hFF;
            15'd1957: data <= 8'hFF;
            15'd1958: data <= 8'hFF;
            15'd1959: data <= 8'hFF;
            15'd1960: data <= 8'hFF;
            15'd1961: data <= 8'hFF;
            15'd1962: data <= 8'hFE;
            15'd1963: data <= 8'h07;
            15'd1964: data <= 8'hFF;
            15'd1965: data <= 8'hFF;
            15'd1966: data <= 8'hE0;
            15'd1967: data <= 8'h7F;
            15'd1968: data <= 8'hFF;
            15'd1969: data <= 8'hFF;
            15'd1970: data <= 8'hFF;
            15'd1971: data <= 8'hFF;
            15'd1972: data <= 8'hFF;
            15'd1973: data <= 8'hFF;
            15'd1974: data <= 8'hFF;
            15'd1975: data <= 8'h80;
            15'd1976: data <= 8'h00;
            15'd1977: data <= 8'h00;
            15'd1978: data <= 8'h00;
            15'd1979: data <= 8'h00;
            15'd1980: data <= 8'h00;
            15'd1981: data <= 8'h00;
            15'd1982: data <= 8'h00;
            15'd1983: data <= 8'h00;
            15'd1984: data <= 8'h01;
            15'd1985: data <= 8'hFF;
            15'd1986: data <= 8'hFF;
            15'd1987: data <= 8'hFF;
            15'd1988: data <= 8'hFF;
            15'd1989: data <= 8'hFF;
            15'd1990: data <= 8'hFF;
            15'd1991: data <= 8'hFF;
            15'd1992: data <= 8'hFF;
            15'd1993: data <= 8'h1F;
            15'd1994: data <= 8'hFF;
            15'd1995: data <= 8'hFF;
            15'd1996: data <= 8'hF9;
            15'd1997: data <= 8'hFF;
            15'd1998: data <= 8'hFF;
            15'd1999: data <= 8'hFF;
            15'd2000: data <= 8'hFF;
            15'd2001: data <= 8'hFF;
            15'd2002: data <= 8'hFF;
            15'd2003: data <= 8'hFF;
            15'd2004: data <= 8'hFF;
            15'd2005: data <= 8'h80;
            15'd2006: data <= 8'h00;
            15'd2007: data <= 8'h00;
            15'd2008: data <= 8'h00;
            15'd2009: data <= 8'h00;
            15'd2010: data <= 8'h00;
            15'd2011: data <= 8'h00;
            15'd2012: data <= 8'h00;
            15'd2013: data <= 8'h00;
            15'd2014: data <= 8'h01;
            15'd2015: data <= 8'hFF;
            15'd2016: data <= 8'hFF;
            15'd2017: data <= 8'hFF;
            15'd2018: data <= 8'hFF;
            15'd2019: data <= 8'hFF;
            15'd2020: data <= 8'hFF;
            15'd2021: data <= 8'hFF;
            15'd2022: data <= 8'hFF;
            15'd2023: data <= 8'hFF;
            15'd2024: data <= 8'hFF;
            15'd2025: data <= 8'hFF;
            15'd2026: data <= 8'hFF;
            15'd2027: data <= 8'hFF;
            15'd2028: data <= 8'hFF;
            15'd2029: data <= 8'hFF;
            15'd2030: data <= 8'hFF;
            15'd2031: data <= 8'hFF;
            15'd2032: data <= 8'hFF;
            15'd2033: data <= 8'hFF;
            15'd2034: data <= 8'hFF;
            15'd2035: data <= 8'h80;
            15'd2036: data <= 8'h00;
            15'd2037: data <= 8'h00;
            15'd2038: data <= 8'h00;
            15'd2039: data <= 8'h00;
            15'd2040: data <= 8'h00;
            15'd2041: data <= 8'h00;
            15'd2042: data <= 8'h00;
            15'd2043: data <= 8'h00;
            15'd2044: data <= 8'h01;
            15'd2045: data <= 8'hFF;
            15'd2046: data <= 8'hFF;
            15'd2047: data <= 8'hFF;
            15'd2048: data <= 8'hFF;
            15'd2049: data <= 8'hFF;
            15'd2050: data <= 8'hFF;
            15'd2051: data <= 8'hFF;
            15'd2052: data <= 8'hFF;
            15'd2053: data <= 8'hFF;
            15'd2054: data <= 8'hFF;
            15'd2055: data <= 8'hFF;
            15'd2056: data <= 8'hFF;
            15'd2057: data <= 8'hFF;
            15'd2058: data <= 8'hFF;
            15'd2059: data <= 8'hFF;
            15'd2060: data <= 8'hFF;
            15'd2061: data <= 8'hFF;
            15'd2062: data <= 8'hFF;
            15'd2063: data <= 8'hFF;
            15'd2064: data <= 8'hFF;
            15'd2065: data <= 8'h80;
            15'd2066: data <= 8'h00;
            15'd2067: data <= 8'h00;
            15'd2068: data <= 8'h00;
            15'd2069: data <= 8'h00;
            15'd2070: data <= 8'h00;
            15'd2071: data <= 8'h00;
            15'd2072: data <= 8'h00;
            15'd2073: data <= 8'h00;
            15'd2074: data <= 8'h01;
            15'd2075: data <= 8'hFF;
            15'd2076: data <= 8'hFF;
            15'd2077: data <= 8'hFF;
            15'd2078: data <= 8'hFF;
            15'd2079: data <= 8'hFF;
            15'd2080: data <= 8'hFF;
            15'd2081: data <= 8'hFF;
            15'd2082: data <= 8'hFF;
            15'd2083: data <= 8'hFF;
            15'd2084: data <= 8'hFF;
            15'd2085: data <= 8'hFF;
            15'd2086: data <= 8'hFF;
            15'd2087: data <= 8'hFF;
            15'd2088: data <= 8'hFF;
            15'd2089: data <= 8'hFF;
            15'd2090: data <= 8'hFF;
            15'd2091: data <= 8'hFF;
            15'd2092: data <= 8'hFF;
            15'd2093: data <= 8'hFF;
            15'd2094: data <= 8'hFF;
            15'd2095: data <= 8'h80;
            15'd2096: data <= 8'h00;
            15'd2097: data <= 8'h00;
            15'd2098: data <= 8'h00;
            15'd2099: data <= 8'h00;
            15'd2100: data <= 8'h00;
            15'd2101: data <= 8'h00;
            15'd2102: data <= 8'h00;
            15'd2103: data <= 8'h00;
            15'd2104: data <= 8'h01;
            15'd2105: data <= 8'hFF;
            15'd2106: data <= 8'hFF;
            15'd2107: data <= 8'hFF;
            15'd2108: data <= 8'hFF;
            15'd2109: data <= 8'hFF;
            15'd2110: data <= 8'hFF;
            15'd2111: data <= 8'hFF;
            15'd2112: data <= 8'hFF;
            15'd2113: data <= 8'hFF;
            15'd2114: data <= 8'hFF;
            15'd2115: data <= 8'hFF;
            15'd2116: data <= 8'hFF;
            15'd2117: data <= 8'hFF;
            15'd2118: data <= 8'hFF;
            15'd2119: data <= 8'hFF;
            15'd2120: data <= 8'hFF;
            15'd2121: data <= 8'hFF;
            15'd2122: data <= 8'hFF;
            15'd2123: data <= 8'hFF;
            15'd2124: data <= 8'hFF;
            15'd2125: data <= 8'h80;
            15'd2126: data <= 8'h00;
            15'd2127: data <= 8'h00;
            15'd2128: data <= 8'h00;
            15'd2129: data <= 8'h00;
            15'd2130: data <= 8'h00;
            15'd2131: data <= 8'h00;
            15'd2132: data <= 8'h00;
            15'd2133: data <= 8'h00;
            15'd2134: data <= 8'h01;
            15'd2135: data <= 8'hFF;
            15'd2136: data <= 8'hFF;
            15'd2137: data <= 8'hFF;
            15'd2138: data <= 8'hFF;
            15'd2139: data <= 8'hFF;
            15'd2140: data <= 8'hFF;
            15'd2141: data <= 8'hFE;
            15'd2142: data <= 8'h7F;
            15'd2143: data <= 8'hFF;
            15'd2144: data <= 8'hFF;
            15'd2145: data <= 8'hFF;
            15'd2146: data <= 8'hFF;
            15'd2147: data <= 8'hFF;
            15'd2148: data <= 8'hF1;
            15'd2149: data <= 8'hF1;
            15'd2150: data <= 8'hFF;
            15'd2151: data <= 8'hFF;
            15'd2152: data <= 8'hFF;
            15'd2153: data <= 8'hFF;
            15'd2154: data <= 8'hFF;
            15'd2155: data <= 8'h80;
            15'd2156: data <= 8'h00;
            15'd2157: data <= 8'h00;
            15'd2158: data <= 8'h00;
            15'd2159: data <= 8'h00;
            15'd2160: data <= 8'h00;
            15'd2161: data <= 8'h00;
            15'd2162: data <= 8'h00;
            15'd2163: data <= 8'h00;
            15'd2164: data <= 8'h01;
            15'd2165: data <= 8'hFF;
            15'd2166: data <= 8'hFF;
            15'd2167: data <= 8'hFF;
            15'd2168: data <= 8'hFF;
            15'd2169: data <= 8'hFF;
            15'd2170: data <= 8'hFF;
            15'd2171: data <= 8'h9C;
            15'd2172: data <= 8'h3F;
            15'd2173: data <= 8'hFF;
            15'd2174: data <= 8'hFF;
            15'd2175: data <= 8'hFF;
            15'd2176: data <= 8'hFF;
            15'd2177: data <= 8'hFF;
            15'd2178: data <= 8'hF0;
            15'd2179: data <= 8'hF1;
            15'd2180: data <= 8'hFF;
            15'd2181: data <= 8'hFF;
            15'd2182: data <= 8'hFF;
            15'd2183: data <= 8'hFF;
            15'd2184: data <= 8'hFF;
            15'd2185: data <= 8'h80;
            15'd2186: data <= 8'h00;
            15'd2187: data <= 8'h00;
            15'd2188: data <= 8'h00;
            15'd2189: data <= 8'h00;
            15'd2190: data <= 8'h00;
            15'd2191: data <= 8'h00;
            15'd2192: data <= 8'h00;
            15'd2193: data <= 8'h00;
            15'd2194: data <= 8'h01;
            15'd2195: data <= 8'hFF;
            15'd2196: data <= 8'hFF;
            15'd2197: data <= 8'hFF;
            15'd2198: data <= 8'hFF;
            15'd2199: data <= 8'hFF;
            15'd2200: data <= 8'hFF;
            15'd2201: data <= 8'h0C;
            15'd2202: data <= 8'h1F;
            15'd2203: data <= 8'hFF;
            15'd2204: data <= 8'hFE;
            15'd2205: data <= 8'h07;
            15'd2206: data <= 8'hFF;
            15'd2207: data <= 8'hFF;
            15'd2208: data <= 8'hE1;
            15'd2209: data <= 8'hE1;
            15'd2210: data <= 8'hFF;
            15'd2211: data <= 8'hFF;
            15'd2212: data <= 8'hFF;
            15'd2213: data <= 8'hFF;
            15'd2214: data <= 8'hFF;
            15'd2215: data <= 8'h80;
            15'd2216: data <= 8'h00;
            15'd2217: data <= 8'h00;
            15'd2218: data <= 8'h00;
            15'd2219: data <= 8'h00;
            15'd2220: data <= 8'h00;
            15'd2221: data <= 8'h00;
            15'd2222: data <= 8'h00;
            15'd2223: data <= 8'h00;
            15'd2224: data <= 8'h01;
            15'd2225: data <= 8'hFF;
            15'd2226: data <= 8'hFF;
            15'd2227: data <= 8'hFF;
            15'd2228: data <= 8'hFF;
            15'd2229: data <= 8'hFF;
            15'd2230: data <= 8'hFE;
            15'd2231: data <= 8'h0C;
            15'd2232: data <= 8'h3F;
            15'd2233: data <= 8'hFF;
            15'd2234: data <= 8'hF8;
            15'd2235: data <= 8'h01;
            15'd2236: data <= 8'hFF;
            15'd2237: data <= 8'hFF;
            15'd2238: data <= 8'hE1;
            15'd2239: data <= 8'hE1;
            15'd2240: data <= 8'hFF;
            15'd2241: data <= 8'hFF;
            15'd2242: data <= 8'hFF;
            15'd2243: data <= 8'hFF;
            15'd2244: data <= 8'hFF;
            15'd2245: data <= 8'h80;
            15'd2246: data <= 8'h00;
            15'd2247: data <= 8'h00;
            15'd2248: data <= 8'h00;
            15'd2249: data <= 8'h00;
            15'd2250: data <= 8'h00;
            15'd2251: data <= 8'h00;
            15'd2252: data <= 8'h00;
            15'd2253: data <= 8'h00;
            15'd2254: data <= 8'h01;
            15'd2255: data <= 8'hFF;
            15'd2256: data <= 8'hFF;
            15'd2257: data <= 8'hFF;
            15'd2258: data <= 8'hFF;
            15'd2259: data <= 8'hFF;
            15'd2260: data <= 8'hFE;
            15'd2261: data <= 8'h1C;
            15'd2262: data <= 8'h3F;
            15'd2263: data <= 8'hFF;
            15'd2264: data <= 8'hF0;
            15'd2265: data <= 8'h00;
            15'd2266: data <= 8'hFF;
            15'd2267: data <= 8'hFF;
            15'd2268: data <= 8'hF1;
            15'd2269: data <= 8'hF1;
            15'd2270: data <= 8'hFF;
            15'd2271: data <= 8'hFF;
            15'd2272: data <= 8'hFF;
            15'd2273: data <= 8'hFF;
            15'd2274: data <= 8'hFF;
            15'd2275: data <= 8'h80;
            15'd2276: data <= 8'h00;
            15'd2277: data <= 8'h00;
            15'd2278: data <= 8'h00;
            15'd2279: data <= 8'h00;
            15'd2280: data <= 8'h00;
            15'd2281: data <= 8'h00;
            15'd2282: data <= 8'h00;
            15'd2283: data <= 8'h00;
            15'd2284: data <= 8'h01;
            15'd2285: data <= 8'hFF;
            15'd2286: data <= 8'hFF;
            15'd2287: data <= 8'hFF;
            15'd2288: data <= 8'hFF;
            15'd2289: data <= 8'hFF;
            15'd2290: data <= 8'hFE;
            15'd2291: data <= 8'h1C;
            15'd2292: data <= 8'h7F;
            15'd2293: data <= 8'hFF;
            15'd2294: data <= 8'hE0;
            15'd2295: data <= 8'h00;
            15'd2296: data <= 8'h7F;
            15'd2297: data <= 8'hFF;
            15'd2298: data <= 8'hF3;
            15'd2299: data <= 8'hF3;
            15'd2300: data <= 8'hFF;
            15'd2301: data <= 8'hFF;
            15'd2302: data <= 8'hFF;
            15'd2303: data <= 8'hFF;
            15'd2304: data <= 8'hFF;
            15'd2305: data <= 8'h80;
            15'd2306: data <= 8'h00;
            15'd2307: data <= 8'h00;
            15'd2308: data <= 8'h00;
            15'd2309: data <= 8'h00;
            15'd2310: data <= 8'h00;
            15'd2311: data <= 8'h00;
            15'd2312: data <= 8'h00;
            15'd2313: data <= 8'h00;
            15'd2314: data <= 8'h01;
            15'd2315: data <= 8'hFF;
            15'd2316: data <= 8'hFF;
            15'd2317: data <= 8'hFF;
            15'd2318: data <= 8'hFF;
            15'd2319: data <= 8'hFF;
            15'd2320: data <= 8'hFF;
            15'd2321: data <= 8'h1C;
            15'd2322: data <= 8'hFF;
            15'd2323: data <= 8'hFF;
            15'd2324: data <= 8'hC0;
            15'd2325: data <= 8'h40;
            15'd2326: data <= 8'h3F;
            15'd2327: data <= 8'hF8;
            15'd2328: data <= 8'hFF;
            15'd2329: data <= 8'hFF;
            15'd2330: data <= 8'hFF;
            15'd2331: data <= 8'hFF;
            15'd2332: data <= 8'hFF;
            15'd2333: data <= 8'hFF;
            15'd2334: data <= 8'hFF;
            15'd2335: data <= 8'h80;
            15'd2336: data <= 8'h00;
            15'd2337: data <= 8'h00;
            15'd2338: data <= 8'h00;
            15'd2339: data <= 8'h00;
            15'd2340: data <= 8'h00;
            15'd2341: data <= 8'h00;
            15'd2342: data <= 8'h00;
            15'd2343: data <= 8'h00;
            15'd2344: data <= 8'h01;
            15'd2345: data <= 8'hFF;
            15'd2346: data <= 8'hFF;
            15'd2347: data <= 8'hFF;
            15'd2348: data <= 8'hFF;
            15'd2349: data <= 8'hFF;
            15'd2350: data <= 8'hFF;
            15'd2351: data <= 8'hBF;
            15'd2352: data <= 8'hFF;
            15'd2353: data <= 8'hFF;
            15'd2354: data <= 8'h81;
            15'd2355: data <= 8'hF0;
            15'd2356: data <= 8'h1F;
            15'd2357: data <= 8'hF8;
            15'd2358: data <= 8'h7F;
            15'd2359: data <= 8'hFF;
            15'd2360: data <= 8'hFF;
            15'd2361: data <= 8'hFF;
            15'd2362: data <= 8'hFF;
            15'd2363: data <= 8'hFF;
            15'd2364: data <= 8'hFF;
            15'd2365: data <= 8'h80;
            15'd2366: data <= 8'h00;
            15'd2367: data <= 8'h00;
            15'd2368: data <= 8'h00;
            15'd2369: data <= 8'h00;
            15'd2370: data <= 8'h00;
            15'd2371: data <= 8'h00;
            15'd2372: data <= 8'h00;
            15'd2373: data <= 8'h00;
            15'd2374: data <= 8'h01;
            15'd2375: data <= 8'hFF;
            15'd2376: data <= 8'hFF;
            15'd2377: data <= 8'hFF;
            15'd2378: data <= 8'hFF;
            15'd2379: data <= 8'hFF;
            15'd2380: data <= 8'hFF;
            15'd2381: data <= 8'hFF;
            15'd2382: data <= 8'hFF;
            15'd2383: data <= 8'hFF;
            15'd2384: data <= 8'h83;
            15'd2385: data <= 8'hFC;
            15'd2386: data <= 8'h1F;
            15'd2387: data <= 8'hF0;
            15'd2388: data <= 8'h7F;
            15'd2389: data <= 8'hFF;
            15'd2390: data <= 8'hFF;
            15'd2391: data <= 8'hFF;
            15'd2392: data <= 8'hFF;
            15'd2393: data <= 8'hFF;
            15'd2394: data <= 8'hFF;
            15'd2395: data <= 8'h80;
            15'd2396: data <= 8'h00;
            15'd2397: data <= 8'h00;
            15'd2398: data <= 8'h00;
            15'd2399: data <= 8'h00;
            15'd2400: data <= 8'h00;
            15'd2401: data <= 8'h00;
            15'd2402: data <= 8'h00;
            15'd2403: data <= 8'h00;
            15'd2404: data <= 8'h01;
            15'd2405: data <= 8'hFF;
            15'd2406: data <= 8'hFF;
            15'd2407: data <= 8'hFF;
            15'd2408: data <= 8'hFF;
            15'd2409: data <= 8'hFF;
            15'd2410: data <= 8'hFF;
            15'd2411: data <= 8'hFF;
            15'd2412: data <= 8'hFF;
            15'd2413: data <= 8'hFF;
            15'd2414: data <= 8'h07;
            15'd2415: data <= 8'hFE;
            15'd2416: data <= 8'h1F;
            15'd2417: data <= 8'hE0;
            15'd2418: data <= 8'hFF;
            15'd2419: data <= 8'hFF;
            15'd2420: data <= 8'hFF;
            15'd2421: data <= 8'hFF;
            15'd2422: data <= 8'hFF;
            15'd2423: data <= 8'hFF;
            15'd2424: data <= 8'hFF;
            15'd2425: data <= 8'h80;
            15'd2426: data <= 8'h00;
            15'd2427: data <= 8'h00;
            15'd2428: data <= 8'h00;
            15'd2429: data <= 8'h00;
            15'd2430: data <= 8'h00;
            15'd2431: data <= 8'h00;
            15'd2432: data <= 8'h00;
            15'd2433: data <= 8'h00;
            15'd2434: data <= 8'h01;
            15'd2435: data <= 8'hFF;
            15'd2436: data <= 8'hFF;
            15'd2437: data <= 8'hFF;
            15'd2438: data <= 8'hFF;
            15'd2439: data <= 8'hFF;
            15'd2440: data <= 8'hFF;
            15'd2441: data <= 8'hFF;
            15'd2442: data <= 8'hFF;
            15'd2443: data <= 8'hFF;
            15'd2444: data <= 8'h0F;
            15'd2445: data <= 8'hFF;
            15'd2446: data <= 8'hFF;
            15'd2447: data <= 8'hE0;
            15'd2448: data <= 8'hFF;
            15'd2449: data <= 8'hFF;
            15'd2450: data <= 8'hFF;
            15'd2451: data <= 8'hFF;
            15'd2452: data <= 8'hFF;
            15'd2453: data <= 8'hFF;
            15'd2454: data <= 8'hFF;
            15'd2455: data <= 8'h80;
            15'd2456: data <= 8'h00;
            15'd2457: data <= 8'h00;
            15'd2458: data <= 8'h00;
            15'd2459: data <= 8'h00;
            15'd2460: data <= 8'h00;
            15'd2461: data <= 8'h00;
            15'd2462: data <= 8'h00;
            15'd2463: data <= 8'h00;
            15'd2464: data <= 8'h01;
            15'd2465: data <= 8'hFF;
            15'd2466: data <= 8'hFF;
            15'd2467: data <= 8'hFF;
            15'd2468: data <= 8'hFF;
            15'd2469: data <= 8'hFF;
            15'd2470: data <= 8'hFF;
            15'd2471: data <= 8'hFF;
            15'd2472: data <= 8'hFF;
            15'd2473: data <= 8'hFF;
            15'd2474: data <= 8'h9F;
            15'd2475: data <= 8'hFF;
            15'd2476: data <= 8'hFF;
            15'd2477: data <= 8'hC1;
            15'd2478: data <= 8'hFF;
            15'd2479: data <= 8'hFF;
            15'd2480: data <= 8'hFF;
            15'd2481: data <= 8'hFF;
            15'd2482: data <= 8'hFF;
            15'd2483: data <= 8'hFF;
            15'd2484: data <= 8'hFF;
            15'd2485: data <= 8'h80;
            15'd2486: data <= 8'h00;
            15'd2487: data <= 8'h00;
            15'd2488: data <= 8'h00;
            15'd2489: data <= 8'h00;
            15'd2490: data <= 8'h00;
            15'd2491: data <= 8'h00;
            15'd2492: data <= 8'h00;
            15'd2493: data <= 8'h00;
            15'd2494: data <= 8'h01;
            15'd2495: data <= 8'hFF;
            15'd2496: data <= 8'hFF;
            15'd2497: data <= 8'hFF;
            15'd2498: data <= 8'hFF;
            15'd2499: data <= 8'hFF;
            15'd2500: data <= 8'hFF;
            15'd2501: data <= 8'hFF;
            15'd2502: data <= 8'hFF;
            15'd2503: data <= 8'hFF;
            15'd2504: data <= 8'hFF;
            15'd2505: data <= 8'hFF;
            15'd2506: data <= 8'hFF;
            15'd2507: data <= 8'hC3;
            15'd2508: data <= 8'hFF;
            15'd2509: data <= 8'hFF;
            15'd2510: data <= 8'hFF;
            15'd2511: data <= 8'hFF;
            15'd2512: data <= 8'hFF;
            15'd2513: data <= 8'hFF;
            15'd2514: data <= 8'hFF;
            15'd2515: data <= 8'h80;
            15'd2516: data <= 8'h00;
            15'd2517: data <= 8'h00;
            15'd2518: data <= 8'h00;
            15'd2519: data <= 8'h00;
            15'd2520: data <= 8'h00;
            15'd2521: data <= 8'h00;
            15'd2522: data <= 8'h00;
            15'd2523: data <= 8'h00;
            15'd2524: data <= 8'h01;
            15'd2525: data <= 8'hFF;
            15'd2526: data <= 8'hFF;
            15'd2527: data <= 8'hFF;
            15'd2528: data <= 8'hFF;
            15'd2529: data <= 8'hFF;
            15'd2530: data <= 8'hFF;
            15'd2531: data <= 8'hFF;
            15'd2532: data <= 8'hFF;
            15'd2533: data <= 8'hFF;
            15'd2534: data <= 8'hFF;
            15'd2535: data <= 8'hFF;
            15'd2536: data <= 8'hFF;
            15'd2537: data <= 8'h83;
            15'd2538: data <= 8'hFF;
            15'd2539: data <= 8'hFF;
            15'd2540: data <= 8'hFF;
            15'd2541: data <= 8'hFF;
            15'd2542: data <= 8'hFF;
            15'd2543: data <= 8'hFF;
            15'd2544: data <= 8'hFF;
            15'd2545: data <= 8'h80;
            15'd2546: data <= 8'h00;
            15'd2547: data <= 8'h00;
            15'd2548: data <= 8'h00;
            15'd2549: data <= 8'h00;
            15'd2550: data <= 8'h00;
            15'd2551: data <= 8'h00;
            15'd2552: data <= 8'h00;
            15'd2553: data <= 8'h00;
            15'd2554: data <= 8'h01;
            15'd2555: data <= 8'hFF;
            15'd2556: data <= 8'hFF;
            15'd2557: data <= 8'hFF;
            15'd2558: data <= 8'hFF;
            15'd2559: data <= 8'hFF;
            15'd2560: data <= 8'hFF;
            15'd2561: data <= 8'hFF;
            15'd2562: data <= 8'hFF;
            15'd2563: data <= 8'hFF;
            15'd2564: data <= 8'hFF;
            15'd2565: data <= 8'hFF;
            15'd2566: data <= 8'hFF;
            15'd2567: data <= 8'h87;
            15'd2568: data <= 8'hFF;
            15'd2569: data <= 8'h1F;
            15'd2570: data <= 8'hFF;
            15'd2571: data <= 8'hFF;
            15'd2572: data <= 8'hFF;
            15'd2573: data <= 8'hFF;
            15'd2574: data <= 8'hFF;
            15'd2575: data <= 8'h80;
            15'd2576: data <= 8'h00;
            15'd2577: data <= 8'h00;
            15'd2578: data <= 8'h00;
            15'd2579: data <= 8'h00;
            15'd2580: data <= 8'h00;
            15'd2581: data <= 8'h00;
            15'd2582: data <= 8'h00;
            15'd2583: data <= 8'h00;
            15'd2584: data <= 8'h01;
            15'd2585: data <= 8'hFF;
            15'd2586: data <= 8'hFF;
            15'd2587: data <= 8'hFF;
            15'd2588: data <= 8'hFF;
            15'd2589: data <= 8'hFF;
            15'd2590: data <= 8'hFF;
            15'd2591: data <= 8'hFF;
            15'd2592: data <= 8'hFF;
            15'd2593: data <= 8'hFF;
            15'd2594: data <= 8'hFF;
            15'd2595: data <= 8'hFF;
            15'd2596: data <= 8'hFF;
            15'd2597: data <= 8'h07;
            15'd2598: data <= 8'hFE;
            15'd2599: data <= 8'h1F;
            15'd2600: data <= 8'hFF;
            15'd2601: data <= 8'hFF;
            15'd2602: data <= 8'hFF;
            15'd2603: data <= 8'hFF;
            15'd2604: data <= 8'hFF;
            15'd2605: data <= 8'h80;
            15'd2606: data <= 8'h00;
            15'd2607: data <= 8'h00;
            15'd2608: data <= 8'h00;
            15'd2609: data <= 8'h00;
            15'd2610: data <= 8'h00;
            15'd2611: data <= 8'h00;
            15'd2612: data <= 8'h00;
            15'd2613: data <= 8'h00;
            15'd2614: data <= 8'h01;
            15'd2615: data <= 8'hFF;
            15'd2616: data <= 8'hFF;
            15'd2617: data <= 8'hFF;
            15'd2618: data <= 8'hFF;
            15'd2619: data <= 8'hFF;
            15'd2620: data <= 8'hFF;
            15'd2621: data <= 8'hFF;
            15'd2622: data <= 8'hFF;
            15'd2623: data <= 8'hFF;
            15'd2624: data <= 8'hFF;
            15'd2625: data <= 8'hFF;
            15'd2626: data <= 8'hFE;
            15'd2627: data <= 8'h0F;
            15'd2628: data <= 8'hFC;
            15'd2629: data <= 8'h1F;
            15'd2630: data <= 8'hFF;
            15'd2631: data <= 8'hFF;
            15'd2632: data <= 8'hFF;
            15'd2633: data <= 8'hFF;
            15'd2634: data <= 8'hFF;
            15'd2635: data <= 8'h80;
            15'd2636: data <= 8'h00;
            15'd2637: data <= 8'h00;
            15'd2638: data <= 8'h00;
            15'd2639: data <= 8'h00;
            15'd2640: data <= 8'h00;
            15'd2641: data <= 8'h00;
            15'd2642: data <= 8'h00;
            15'd2643: data <= 8'h00;
            15'd2644: data <= 8'h01;
            15'd2645: data <= 8'hFF;
            15'd2646: data <= 8'hFF;
            15'd2647: data <= 8'hFF;
            15'd2648: data <= 8'hFF;
            15'd2649: data <= 8'hFF;
            15'd2650: data <= 8'hFF;
            15'd2651: data <= 8'hFF;
            15'd2652: data <= 8'hFF;
            15'd2653: data <= 8'hFF;
            15'd2654: data <= 8'hFF;
            15'd2655: data <= 8'hFF;
            15'd2656: data <= 8'hFE;
            15'd2657: data <= 8'h0F;
            15'd2658: data <= 8'hF8;
            15'd2659: data <= 8'h3F;
            15'd2660: data <= 8'hFF;
            15'd2661: data <= 8'hFF;
            15'd2662: data <= 8'hFF;
            15'd2663: data <= 8'hFF;
            15'd2664: data <= 8'hFF;
            15'd2665: data <= 8'h80;
            15'd2666: data <= 8'h00;
            15'd2667: data <= 8'h00;
            15'd2668: data <= 8'h00;
            15'd2669: data <= 8'h00;
            15'd2670: data <= 8'h00;
            15'd2671: data <= 8'h00;
            15'd2672: data <= 8'h00;
            15'd2673: data <= 8'h00;
            15'd2674: data <= 8'h01;
            15'd2675: data <= 8'hFF;
            15'd2676: data <= 8'hFF;
            15'd2677: data <= 8'hFF;
            15'd2678: data <= 8'hFF;
            15'd2679: data <= 8'hFF;
            15'd2680: data <= 8'hFF;
            15'd2681: data <= 8'hFF;
            15'd2682: data <= 8'hFF;
            15'd2683: data <= 8'hFF;
            15'd2684: data <= 8'hFF;
            15'd2685: data <= 8'hFF;
            15'd2686: data <= 8'hFE;
            15'd2687: data <= 8'h1F;
            15'd2688: data <= 8'hF8;
            15'd2689: data <= 8'h3F;
            15'd2690: data <= 8'hFF;
            15'd2691: data <= 8'hFF;
            15'd2692: data <= 8'hFF;
            15'd2693: data <= 8'hFF;
            15'd2694: data <= 8'hFF;
            15'd2695: data <= 8'h80;
            15'd2696: data <= 8'h00;
            15'd2697: data <= 8'h00;
            15'd2698: data <= 8'h00;
            15'd2699: data <= 8'h00;
            15'd2700: data <= 8'h00;
            15'd2701: data <= 8'h00;
            15'd2702: data <= 8'h00;
            15'd2703: data <= 8'h00;
            15'd2704: data <= 8'h01;
            15'd2705: data <= 8'hFF;
            15'd2706: data <= 8'hFF;
            15'd2707: data <= 8'hFF;
            15'd2708: data <= 8'hFF;
            15'd2709: data <= 8'hFF;
            15'd2710: data <= 8'hFF;
            15'd2711: data <= 8'hFF;
            15'd2712: data <= 8'hFF;
            15'd2713: data <= 8'hFF;
            15'd2714: data <= 8'hFF;
            15'd2715: data <= 8'hFF;
            15'd2716: data <= 8'hFC;
            15'd2717: data <= 8'h1F;
            15'd2718: data <= 8'hF0;
            15'd2719: data <= 8'h7F;
            15'd2720: data <= 8'hFF;
            15'd2721: data <= 8'hFF;
            15'd2722: data <= 8'hFF;
            15'd2723: data <= 8'hFF;
            15'd2724: data <= 8'hFF;
            15'd2725: data <= 8'h80;
            15'd2726: data <= 8'h00;
            15'd2727: data <= 8'h00;
            15'd2728: data <= 8'h00;
            15'd2729: data <= 8'h00;
            15'd2730: data <= 8'h00;
            15'd2731: data <= 8'h00;
            15'd2732: data <= 8'h00;
            15'd2733: data <= 8'h00;
            15'd2734: data <= 8'h01;
            15'd2735: data <= 8'hFF;
            15'd2736: data <= 8'hFF;
            15'd2737: data <= 8'hFF;
            15'd2738: data <= 8'hFF;
            15'd2739: data <= 8'hFF;
            15'd2740: data <= 8'hFF;
            15'd2741: data <= 8'hFF;
            15'd2742: data <= 8'hFF;
            15'd2743: data <= 8'hFF;
            15'd2744: data <= 8'hFF;
            15'd2745: data <= 8'hFF;
            15'd2746: data <= 8'hFC;
            15'd2747: data <= 8'h3F;
            15'd2748: data <= 8'hE0;
            15'd2749: data <= 8'hFF;
            15'd2750: data <= 8'hFF;
            15'd2751: data <= 8'hFF;
            15'd2752: data <= 8'hFF;
            15'd2753: data <= 8'hFF;
            15'd2754: data <= 8'hFF;
            15'd2755: data <= 8'h80;
            15'd2756: data <= 8'h00;
            15'd2757: data <= 8'h00;
            15'd2758: data <= 8'h00;
            15'd2759: data <= 8'h00;
            15'd2760: data <= 8'h00;
            15'd2761: data <= 8'h00;
            15'd2762: data <= 8'h00;
            15'd2763: data <= 8'h00;
            15'd2764: data <= 8'h01;
            15'd2765: data <= 8'hFF;
            15'd2766: data <= 8'hFF;
            15'd2767: data <= 8'hFF;
            15'd2768: data <= 8'hFF;
            15'd2769: data <= 8'hFF;
            15'd2770: data <= 8'hFF;
            15'd2771: data <= 8'hFF;
            15'd2772: data <= 8'hFF;
            15'd2773: data <= 8'hFF;
            15'd2774: data <= 8'hFF;
            15'd2775: data <= 8'hFF;
            15'd2776: data <= 8'hFC;
            15'd2777: data <= 8'h3F;
            15'd2778: data <= 8'hC0;
            15'd2779: data <= 8'hFF;
            15'd2780: data <= 8'hFF;
            15'd2781: data <= 8'hFF;
            15'd2782: data <= 8'hFF;
            15'd2783: data <= 8'hFF;
            15'd2784: data <= 8'hFF;
            15'd2785: data <= 8'h80;
            15'd2786: data <= 8'h00;
            15'd2787: data <= 8'h00;
            15'd2788: data <= 8'h00;
            15'd2789: data <= 8'h00;
            15'd2790: data <= 8'h00;
            15'd2791: data <= 8'h00;
            15'd2792: data <= 8'h00;
            15'd2793: data <= 8'h00;
            15'd2794: data <= 8'h01;
            15'd2795: data <= 8'hFF;
            15'd2796: data <= 8'hFF;
            15'd2797: data <= 8'hFF;
            15'd2798: data <= 8'hFF;
            15'd2799: data <= 8'hFF;
            15'd2800: data <= 8'hFF;
            15'd2801: data <= 8'hFF;
            15'd2802: data <= 8'hFF;
            15'd2803: data <= 8'hFF;
            15'd2804: data <= 8'hFF;
            15'd2805: data <= 8'hFF;
            15'd2806: data <= 8'hF8;
            15'd2807: data <= 8'h7F;
            15'd2808: data <= 8'h81;
            15'd2809: data <= 8'hFF;
            15'd2810: data <= 8'hFF;
            15'd2811: data <= 8'hFF;
            15'd2812: data <= 8'hFF;
            15'd2813: data <= 8'hFF;
            15'd2814: data <= 8'hFF;
            15'd2815: data <= 8'h80;
            15'd2816: data <= 8'h00;
            15'd2817: data <= 8'h00;
            15'd2818: data <= 8'h00;
            15'd2819: data <= 8'h00;
            15'd2820: data <= 8'h00;
            15'd2821: data <= 8'h00;
            15'd2822: data <= 8'h00;
            15'd2823: data <= 8'h00;
            15'd2824: data <= 8'h01;
            15'd2825: data <= 8'hFF;
            15'd2826: data <= 8'hFF;
            15'd2827: data <= 8'hFF;
            15'd2828: data <= 8'hFF;
            15'd2829: data <= 8'hFF;
            15'd2830: data <= 8'hFF;
            15'd2831: data <= 8'hFF;
            15'd2832: data <= 8'hFF;
            15'd2833: data <= 8'hFF;
            15'd2834: data <= 8'hFF;
            15'd2835: data <= 8'hFF;
            15'd2836: data <= 8'hF8;
            15'd2837: data <= 8'h7F;
            15'd2838: data <= 8'h03;
            15'd2839: data <= 8'hFF;
            15'd2840: data <= 8'hFF;
            15'd2841: data <= 8'hFF;
            15'd2842: data <= 8'hFF;
            15'd2843: data <= 8'hFF;
            15'd2844: data <= 8'hFF;
            15'd2845: data <= 8'h80;
            15'd2846: data <= 8'h00;
            15'd2847: data <= 8'h00;
            15'd2848: data <= 8'h00;
            15'd2849: data <= 8'h00;
            15'd2850: data <= 8'h00;
            15'd2851: data <= 8'h00;
            15'd2852: data <= 8'h00;
            15'd2853: data <= 8'h00;
            15'd2854: data <= 8'h01;
            15'd2855: data <= 8'hFF;
            15'd2856: data <= 8'hFF;
            15'd2857: data <= 8'hFF;
            15'd2858: data <= 8'hFF;
            15'd2859: data <= 8'hFF;
            15'd2860: data <= 8'hFF;
            15'd2861: data <= 8'hFF;
            15'd2862: data <= 8'hFF;
            15'd2863: data <= 8'hFF;
            15'd2864: data <= 8'hFF;
            15'd2865: data <= 8'hFF;
            15'd2866: data <= 8'hF8;
            15'd2867: data <= 8'h7E;
            15'd2868: data <= 8'h07;
            15'd2869: data <= 8'hFF;
            15'd2870: data <= 8'hFF;
            15'd2871: data <= 8'hFF;
            15'd2872: data <= 8'hFF;
            15'd2873: data <= 8'hFF;
            15'd2874: data <= 8'hFF;
            15'd2875: data <= 8'h80;
            15'd2876: data <= 8'h00;
            15'd2877: data <= 8'h00;
            15'd2878: data <= 8'h00;
            15'd2879: data <= 8'h00;
            15'd2880: data <= 8'h00;
            15'd2881: data <= 8'h00;
            15'd2882: data <= 8'h00;
            15'd2883: data <= 8'h00;
            15'd2884: data <= 8'h01;
            15'd2885: data <= 8'hFF;
            15'd2886: data <= 8'hFF;
            15'd2887: data <= 8'hFF;
            15'd2888: data <= 8'hFF;
            15'd2889: data <= 8'hFF;
            15'd2890: data <= 8'hFF;
            15'd2891: data <= 8'hFF;
            15'd2892: data <= 8'hFF;
            15'd2893: data <= 8'hFF;
            15'd2894: data <= 8'hFF;
            15'd2895: data <= 8'hFF;
            15'd2896: data <= 8'hF8;
            15'd2897: data <= 8'h7C;
            15'd2898: data <= 8'h0F;
            15'd2899: data <= 8'hFF;
            15'd2900: data <= 8'hFF;
            15'd2901: data <= 8'hFF;
            15'd2902: data <= 8'hFF;
            15'd2903: data <= 8'hFF;
            15'd2904: data <= 8'hFF;
            15'd2905: data <= 8'h80;
            15'd2906: data <= 8'h00;
            15'd2907: data <= 8'h00;
            15'd2908: data <= 8'h00;
            15'd2909: data <= 8'h00;
            15'd2910: data <= 8'h00;
            15'd2911: data <= 8'h00;
            15'd2912: data <= 8'h00;
            15'd2913: data <= 8'h00;
            15'd2914: data <= 8'h01;
            15'd2915: data <= 8'hFF;
            15'd2916: data <= 8'hFF;
            15'd2917: data <= 8'hFF;
            15'd2918: data <= 8'hFF;
            15'd2919: data <= 8'hFF;
            15'd2920: data <= 8'hFF;
            15'd2921: data <= 8'hFF;
            15'd2922: data <= 8'hFF;
            15'd2923: data <= 8'hFF;
            15'd2924: data <= 8'hFF;
            15'd2925: data <= 8'hFF;
            15'd2926: data <= 8'hF8;
            15'd2927: data <= 8'h70;
            15'd2928: data <= 8'h1F;
            15'd2929: data <= 8'hFF;
            15'd2930: data <= 8'hFF;
            15'd2931: data <= 8'hFF;
            15'd2932: data <= 8'hFF;
            15'd2933: data <= 8'hFF;
            15'd2934: data <= 8'hFF;
            15'd2935: data <= 8'h80;
            15'd2936: data <= 8'h00;
            15'd2937: data <= 8'h00;
            15'd2938: data <= 8'h00;
            15'd2939: data <= 8'h00;
            15'd2940: data <= 8'h00;
            15'd2941: data <= 8'h00;
            15'd2942: data <= 8'h00;
            15'd2943: data <= 8'h00;
            15'd2944: data <= 8'h01;
            15'd2945: data <= 8'hFF;
            15'd2946: data <= 8'hFF;
            15'd2947: data <= 8'hFF;
            15'd2948: data <= 8'hFF;
            15'd2949: data <= 8'hFF;
            15'd2950: data <= 8'hFF;
            15'd2951: data <= 8'hFF;
            15'd2952: data <= 8'hFF;
            15'd2953: data <= 8'hFF;
            15'd2954: data <= 8'hFF;
            15'd2955: data <= 8'hFF;
            15'd2956: data <= 8'hF8;
            15'd2957: data <= 8'h40;
            15'd2958: data <= 8'h3F;
            15'd2959: data <= 8'hFF;
            15'd2960: data <= 8'hFF;
            15'd2961: data <= 8'hFF;
            15'd2962: data <= 8'hFF;
            15'd2963: data <= 8'hFF;
            15'd2964: data <= 8'hFF;
            15'd2965: data <= 8'h80;
            15'd2966: data <= 8'h00;
            15'd2967: data <= 8'h00;
            15'd2968: data <= 8'h00;
            15'd2969: data <= 8'h00;
            15'd2970: data <= 8'h00;
            15'd2971: data <= 8'h00;
            15'd2972: data <= 8'h00;
            15'd2973: data <= 8'h00;
            15'd2974: data <= 8'h01;
            15'd2975: data <= 8'hFF;
            15'd2976: data <= 8'hFF;
            15'd2977: data <= 8'hFF;
            15'd2978: data <= 8'hFF;
            15'd2979: data <= 8'hFF;
            15'd2980: data <= 8'hFF;
            15'd2981: data <= 8'hFF;
            15'd2982: data <= 8'hFF;
            15'd2983: data <= 8'hFF;
            15'd2984: data <= 8'hFF;
            15'd2985: data <= 8'hFF;
            15'd2986: data <= 8'hF8;
            15'd2987: data <= 8'h00;
            15'd2988: data <= 8'h7F;
            15'd2989: data <= 8'hFF;
            15'd2990: data <= 8'hFF;
            15'd2991: data <= 8'hFF;
            15'd2992: data <= 8'hFF;
            15'd2993: data <= 8'hFF;
            15'd2994: data <= 8'hFF;
            15'd2995: data <= 8'h80;
            15'd2996: data <= 8'h00;
            15'd2997: data <= 8'h00;
            15'd2998: data <= 8'h00;
            15'd2999: data <= 8'h00;
            15'd3000: data <= 8'h00;
            15'd3001: data <= 8'h00;
            15'd3002: data <= 8'h00;
            15'd3003: data <= 8'h00;
            15'd3004: data <= 8'h01;
            15'd3005: data <= 8'hFF;
            15'd3006: data <= 8'hFF;
            15'd3007: data <= 8'hFF;
            15'd3008: data <= 8'hFF;
            15'd3009: data <= 8'hFF;
            15'd3010: data <= 8'hFF;
            15'd3011: data <= 8'hFF;
            15'd3012: data <= 8'hFF;
            15'd3013: data <= 8'hFF;
            15'd3014: data <= 8'hFF;
            15'd3015: data <= 8'hFF;
            15'd3016: data <= 8'hFC;
            15'd3017: data <= 8'h00;
            15'd3018: data <= 8'hFF;
            15'd3019: data <= 8'hFF;
            15'd3020: data <= 8'hFF;
            15'd3021: data <= 8'hFF;
            15'd3022: data <= 8'hFF;
            15'd3023: data <= 8'hFF;
            15'd3024: data <= 8'hFF;
            15'd3025: data <= 8'h80;
            15'd3026: data <= 8'h00;
            15'd3027: data <= 8'h00;
            15'd3028: data <= 8'h00;
            15'd3029: data <= 8'h00;
            15'd3030: data <= 8'h00;
            15'd3031: data <= 8'h00;
            15'd3032: data <= 8'h00;
            15'd3033: data <= 8'h00;
            15'd3034: data <= 8'h01;
            15'd3035: data <= 8'hFF;
            15'd3036: data <= 8'hFF;
            15'd3037: data <= 8'hFF;
            15'd3038: data <= 8'hFF;
            15'd3039: data <= 8'hFF;
            15'd3040: data <= 8'hFF;
            15'd3041: data <= 8'hFF;
            15'd3042: data <= 8'hFF;
            15'd3043: data <= 8'hFF;
            15'd3044: data <= 8'hFF;
            15'd3045: data <= 8'hCF;
            15'd3046: data <= 8'hFC;
            15'd3047: data <= 8'h03;
            15'd3048: data <= 8'hFF;
            15'd3049: data <= 8'hFF;
            15'd3050: data <= 8'hFF;
            15'd3051: data <= 8'hFF;
            15'd3052: data <= 8'hFF;
            15'd3053: data <= 8'hFF;
            15'd3054: data <= 8'hFF;
            15'd3055: data <= 8'h80;
            15'd3056: data <= 8'h00;
            15'd3057: data <= 8'h00;
            15'd3058: data <= 8'h00;
            15'd3059: data <= 8'h00;
            15'd3060: data <= 8'h00;
            15'd3061: data <= 8'h00;
            15'd3062: data <= 8'h00;
            15'd3063: data <= 8'h00;
            15'd3064: data <= 8'h01;
            15'd3065: data <= 8'hFF;
            15'd3066: data <= 8'hFF;
            15'd3067: data <= 8'hFF;
            15'd3068: data <= 8'hFF;
            15'd3069: data <= 8'hFF;
            15'd3070: data <= 8'hFF;
            15'd3071: data <= 8'hFF;
            15'd3072: data <= 8'hFF;
            15'd3073: data <= 8'hFF;
            15'd3074: data <= 8'hFF;
            15'd3075: data <= 8'h8F;
            15'd3076: data <= 8'hFF;
            15'd3077: data <= 8'h0F;
            15'd3078: data <= 8'hFF;
            15'd3079: data <= 8'hFF;
            15'd3080: data <= 8'hFF;
            15'd3081: data <= 8'hFF;
            15'd3082: data <= 8'hFF;
            15'd3083: data <= 8'hFF;
            15'd3084: data <= 8'hFF;
            15'd3085: data <= 8'h80;
            15'd3086: data <= 8'h00;
            15'd3087: data <= 8'h00;
            15'd3088: data <= 8'h00;
            15'd3089: data <= 8'h00;
            15'd3090: data <= 8'h00;
            15'd3091: data <= 8'h00;
            15'd3092: data <= 8'h00;
            15'd3093: data <= 8'h00;
            15'd3094: data <= 8'h01;
            15'd3095: data <= 8'hFF;
            15'd3096: data <= 8'hFF;
            15'd3097: data <= 8'hFF;
            15'd3098: data <= 8'hFF;
            15'd3099: data <= 8'hFF;
            15'd3100: data <= 8'hFF;
            15'd3101: data <= 8'hFF;
            15'd3102: data <= 8'hFF;
            15'd3103: data <= 8'hFF;
            15'd3104: data <= 8'hFF;
            15'd3105: data <= 8'h8F;
            15'd3106: data <= 8'hFF;
            15'd3107: data <= 8'hFF;
            15'd3108: data <= 8'hFF;
            15'd3109: data <= 8'hFF;
            15'd3110: data <= 8'hFF;
            15'd3111: data <= 8'hFF;
            15'd3112: data <= 8'hFF;
            15'd3113: data <= 8'hFF;
            15'd3114: data <= 8'hFF;
            15'd3115: data <= 8'h80;
            15'd3116: data <= 8'h00;
            15'd3117: data <= 8'h00;
            15'd3118: data <= 8'h00;
            15'd3119: data <= 8'h00;
            15'd3120: data <= 8'h00;
            15'd3121: data <= 8'h00;
            15'd3122: data <= 8'h00;
            15'd3123: data <= 8'h00;
            15'd3124: data <= 8'h01;
            15'd3125: data <= 8'hFF;
            15'd3126: data <= 8'hFF;
            15'd3127: data <= 8'hFF;
            15'd3128: data <= 8'hFF;
            15'd3129: data <= 8'hFF;
            15'd3130: data <= 8'hFF;
            15'd3131: data <= 8'hFF;
            15'd3132: data <= 8'hFF;
            15'd3133: data <= 8'hFF;
            15'd3134: data <= 8'hFF;
            15'd3135: data <= 8'h1F;
            15'd3136: data <= 8'h7F;
            15'd3137: data <= 8'hFF;
            15'd3138: data <= 8'hFF;
            15'd3139: data <= 8'hFF;
            15'd3140: data <= 8'hFF;
            15'd3141: data <= 8'hFF;
            15'd3142: data <= 8'hFF;
            15'd3143: data <= 8'hFF;
            15'd3144: data <= 8'hFF;
            15'd3145: data <= 8'h80;
            15'd3146: data <= 8'h00;
            15'd3147: data <= 8'h00;
            15'd3148: data <= 8'h00;
            15'd3149: data <= 8'h00;
            15'd3150: data <= 8'h00;
            15'd3151: data <= 8'h00;
            15'd3152: data <= 8'h00;
            15'd3153: data <= 8'h00;
            15'd3154: data <= 8'h01;
            15'd3155: data <= 8'hFF;
            15'd3156: data <= 8'hFF;
            15'd3157: data <= 8'hFF;
            15'd3158: data <= 8'hFF;
            15'd3159: data <= 8'hFF;
            15'd3160: data <= 8'hFF;
            15'd3161: data <= 8'hFF;
            15'd3162: data <= 8'hFF;
            15'd3163: data <= 8'hFF;
            15'd3164: data <= 8'hFE;
            15'd3165: data <= 8'h1E;
            15'd3166: data <= 8'h3F;
            15'd3167: data <= 8'h9F;
            15'd3168: data <= 8'hFF;
            15'd3169: data <= 8'hFF;
            15'd3170: data <= 8'hFF;
            15'd3171: data <= 8'hFF;
            15'd3172: data <= 8'hFF;
            15'd3173: data <= 8'hFF;
            15'd3174: data <= 8'hFF;
            15'd3175: data <= 8'h80;
            15'd3176: data <= 8'h00;
            15'd3177: data <= 8'h00;
            15'd3178: data <= 8'h00;
            15'd3179: data <= 8'h00;
            15'd3180: data <= 8'h00;
            15'd3181: data <= 8'h00;
            15'd3182: data <= 8'h00;
            15'd3183: data <= 8'h00;
            15'd3184: data <= 8'h01;
            15'd3185: data <= 8'hFF;
            15'd3186: data <= 8'hFF;
            15'd3187: data <= 8'hFF;
            15'd3188: data <= 8'hFF;
            15'd3189: data <= 8'hFF;
            15'd3190: data <= 8'hFF;
            15'd3191: data <= 8'hFF;
            15'd3192: data <= 8'hFF;
            15'd3193: data <= 8'hFF;
            15'd3194: data <= 8'hFE;
            15'd3195: data <= 8'h3C;
            15'd3196: data <= 8'h7F;
            15'd3197: data <= 8'h1F;
            15'd3198: data <= 8'hFF;
            15'd3199: data <= 8'hFF;
            15'd3200: data <= 8'hFF;
            15'd3201: data <= 8'hFF;
            15'd3202: data <= 8'hFF;
            15'd3203: data <= 8'hFF;
            15'd3204: data <= 8'hFF;
            15'd3205: data <= 8'h80;
            15'd3206: data <= 8'h00;
            15'd3207: data <= 8'h00;
            15'd3208: data <= 8'h00;
            15'd3209: data <= 8'h00;
            15'd3210: data <= 8'h00;
            15'd3211: data <= 8'h00;
            15'd3212: data <= 8'h00;
            15'd3213: data <= 8'h00;
            15'd3214: data <= 8'h01;
            15'd3215: data <= 8'hFF;
            15'd3216: data <= 8'hFF;
            15'd3217: data <= 8'hFF;
            15'd3218: data <= 8'hFF;
            15'd3219: data <= 8'hFF;
            15'd3220: data <= 8'hFF;
            15'd3221: data <= 8'hFF;
            15'd3222: data <= 8'hFF;
            15'd3223: data <= 8'hFF;
            15'd3224: data <= 8'hFC;
            15'd3225: data <= 8'h7C;
            15'd3226: data <= 8'h7E;
            15'd3227: data <= 8'h1F;
            15'd3228: data <= 8'hFF;
            15'd3229: data <= 8'hFF;
            15'd3230: data <= 8'hFF;
            15'd3231: data <= 8'hFF;
            15'd3232: data <= 8'hFF;
            15'd3233: data <= 8'hFF;
            15'd3234: data <= 8'hFF;
            15'd3235: data <= 8'h80;
            15'd3236: data <= 8'h00;
            15'd3237: data <= 8'h00;
            15'd3238: data <= 8'h00;
            15'd3239: data <= 8'h00;
            15'd3240: data <= 8'h00;
            15'd3241: data <= 8'h00;
            15'd3242: data <= 8'h00;
            15'd3243: data <= 8'h00;
            15'd3244: data <= 8'h01;
            15'd3245: data <= 8'hFF;
            15'd3246: data <= 8'hFF;
            15'd3247: data <= 8'hFF;
            15'd3248: data <= 8'hFF;
            15'd3249: data <= 8'hFF;
            15'd3250: data <= 8'hFF;
            15'd3251: data <= 8'hFF;
            15'd3252: data <= 8'hFF;
            15'd3253: data <= 8'hFF;
            15'd3254: data <= 8'hFF;
            15'd3255: data <= 8'hF8;
            15'd3256: data <= 8'hFE;
            15'd3257: data <= 8'h3F;
            15'd3258: data <= 8'hFF;
            15'd3259: data <= 8'hFF;
            15'd3260: data <= 8'hFF;
            15'd3261: data <= 8'hFF;
            15'd3262: data <= 8'hFF;
            15'd3263: data <= 8'hFF;
            15'd3264: data <= 8'hFF;
            15'd3265: data <= 8'h80;
            15'd3266: data <= 8'h00;
            15'd3267: data <= 8'h00;
            15'd3268: data <= 8'h00;
            15'd3269: data <= 8'h00;
            15'd3270: data <= 8'h00;
            15'd3271: data <= 8'h00;
            15'd3272: data <= 8'h00;
            15'd3273: data <= 8'h00;
            15'd3274: data <= 8'h01;
            15'd3275: data <= 8'hFF;
            15'd3276: data <= 8'hFF;
            15'd3277: data <= 8'hFF;
            15'd3278: data <= 8'hFF;
            15'd3279: data <= 8'hFF;
            15'd3280: data <= 8'hFF;
            15'd3281: data <= 8'hFF;
            15'd3282: data <= 8'hFF;
            15'd3283: data <= 8'hFF;
            15'd3284: data <= 8'hFF;
            15'd3285: data <= 8'hF1;
            15'd3286: data <= 8'hFC;
            15'd3287: data <= 8'h7F;
            15'd3288: data <= 8'hFF;
            15'd3289: data <= 8'hFF;
            15'd3290: data <= 8'hFF;
            15'd3291: data <= 8'hFF;
            15'd3292: data <= 8'hFF;
            15'd3293: data <= 8'hFF;
            15'd3294: data <= 8'hFF;
            15'd3295: data <= 8'h80;
            15'd3296: data <= 8'h00;
            15'd3297: data <= 8'h00;
            15'd3298: data <= 8'h00;
            15'd3299: data <= 8'h00;
            15'd3300: data <= 8'h00;
            15'd3301: data <= 8'h00;
            15'd3302: data <= 8'h00;
            15'd3303: data <= 8'h00;
            15'd3304: data <= 8'h01;
            15'd3305: data <= 8'hFF;
            15'd3306: data <= 8'hFF;
            15'd3307: data <= 8'hFF;
            15'd3308: data <= 8'hFF;
            15'd3309: data <= 8'hFF;
            15'd3310: data <= 8'hFF;
            15'd3311: data <= 8'hFF;
            15'd3312: data <= 8'hFF;
            15'd3313: data <= 8'hFF;
            15'd3314: data <= 8'hFF;
            15'd3315: data <= 8'hF1;
            15'd3316: data <= 8'hF8;
            15'd3317: data <= 8'hFF;
            15'd3318: data <= 8'hFF;
            15'd3319: data <= 8'hFF;
            15'd3320: data <= 8'hFF;
            15'd3321: data <= 8'hFF;
            15'd3322: data <= 8'hFF;
            15'd3323: data <= 8'hFF;
            15'd3324: data <= 8'hFF;
            15'd3325: data <= 8'h80;
            15'd3326: data <= 8'h00;
            15'd3327: data <= 8'h00;
            15'd3328: data <= 8'h00;
            15'd3329: data <= 8'h00;
            15'd3330: data <= 8'h00;
            15'd3331: data <= 8'h00;
            15'd3332: data <= 8'h00;
            15'd3333: data <= 8'h00;
            15'd3334: data <= 8'h01;
            15'd3335: data <= 8'hFF;
            15'd3336: data <= 8'hFF;
            15'd3337: data <= 8'hFF;
            15'd3338: data <= 8'hFF;
            15'd3339: data <= 8'hFF;
            15'd3340: data <= 8'hFF;
            15'd3341: data <= 8'hFF;
            15'd3342: data <= 8'hFF;
            15'd3343: data <= 8'hFF;
            15'd3344: data <= 8'hFF;
            15'd3345: data <= 8'hE3;
            15'd3346: data <= 8'hF0;
            15'd3347: data <= 8'hFF;
            15'd3348: data <= 8'hFF;
            15'd3349: data <= 8'hFF;
            15'd3350: data <= 8'hFF;
            15'd3351: data <= 8'hFF;
            15'd3352: data <= 8'hFF;
            15'd3353: data <= 8'hFF;
            15'd3354: data <= 8'hFF;
            15'd3355: data <= 8'h80;
            15'd3356: data <= 8'h00;
            15'd3357: data <= 8'h00;
            15'd3358: data <= 8'h00;
            15'd3359: data <= 8'h00;
            15'd3360: data <= 8'h00;
            15'd3361: data <= 8'h00;
            15'd3362: data <= 8'h00;
            15'd3363: data <= 8'h00;
            15'd3364: data <= 8'h01;
            15'd3365: data <= 8'hFF;
            15'd3366: data <= 8'hFF;
            15'd3367: data <= 8'hFF;
            15'd3368: data <= 8'hFF;
            15'd3369: data <= 8'hFF;
            15'd3370: data <= 8'hFF;
            15'd3371: data <= 8'hFF;
            15'd3372: data <= 8'hFF;
            15'd3373: data <= 8'hFF;
            15'd3374: data <= 8'hFF;
            15'd3375: data <= 8'hE7;
            15'd3376: data <= 8'hF1;
            15'd3377: data <= 8'hFF;
            15'd3378: data <= 8'hFF;
            15'd3379: data <= 8'hFF;
            15'd3380: data <= 8'hFF;
            15'd3381: data <= 8'hFF;
            15'd3382: data <= 8'hFF;
            15'd3383: data <= 8'hFF;
            15'd3384: data <= 8'hFF;
            15'd3385: data <= 8'h80;
            15'd3386: data <= 8'h00;
            15'd3387: data <= 8'h00;
            15'd3388: data <= 8'h00;
            15'd3389: data <= 8'h00;
            15'd3390: data <= 8'h00;
            15'd3391: data <= 8'h00;
            15'd3392: data <= 8'h00;
            15'd3393: data <= 8'h00;
            15'd3394: data <= 8'h01;
            15'd3395: data <= 8'hFF;
            15'd3396: data <= 8'hFF;
            15'd3397: data <= 8'hFF;
            15'd3398: data <= 8'hFF;
            15'd3399: data <= 8'hFF;
            15'd3400: data <= 8'hFF;
            15'd3401: data <= 8'hFF;
            15'd3402: data <= 8'hFF;
            15'd3403: data <= 8'hC0;
            15'd3404: data <= 8'hFF;
            15'd3405: data <= 8'hEF;
            15'd3406: data <= 8'hE3;
            15'd3407: data <= 8'hFF;
            15'd3408: data <= 8'hFF;
            15'd3409: data <= 8'hFF;
            15'd3410: data <= 8'hFF;
            15'd3411: data <= 8'hFF;
            15'd3412: data <= 8'hFF;
            15'd3413: data <= 8'hFF;
            15'd3414: data <= 8'hFF;
            15'd3415: data <= 8'h80;
            15'd3416: data <= 8'h00;
            15'd3417: data <= 8'h00;
            15'd3418: data <= 8'h00;
            15'd3419: data <= 8'h00;
            15'd3420: data <= 8'h00;
            15'd3421: data <= 8'h00;
            15'd3422: data <= 8'h00;
            15'd3423: data <= 8'h00;
            15'd3424: data <= 8'h01;
            15'd3425: data <= 8'hFF;
            15'd3426: data <= 8'hFF;
            15'd3427: data <= 8'hFF;
            15'd3428: data <= 8'hFF;
            15'd3429: data <= 8'hFF;
            15'd3430: data <= 8'hFF;
            15'd3431: data <= 8'hFF;
            15'd3432: data <= 8'hE3;
            15'd3433: data <= 8'h80;
            15'd3434: data <= 8'h7F;
            15'd3435: data <= 8'hFF;
            15'd3436: data <= 8'hC3;
            15'd3437: data <= 8'hFF;
            15'd3438: data <= 8'hFF;
            15'd3439: data <= 8'hFF;
            15'd3440: data <= 8'hFF;
            15'd3441: data <= 8'hFF;
            15'd3442: data <= 8'hFF;
            15'd3443: data <= 8'hFF;
            15'd3444: data <= 8'hFF;
            15'd3445: data <= 8'h80;
            15'd3446: data <= 8'h00;
            15'd3447: data <= 8'h00;
            15'd3448: data <= 8'h00;
            15'd3449: data <= 8'h00;
            15'd3450: data <= 8'h00;
            15'd3451: data <= 8'h00;
            15'd3452: data <= 8'h00;
            15'd3453: data <= 8'h00;
            15'd3454: data <= 8'h01;
            15'd3455: data <= 8'hFF;
            15'd3456: data <= 8'hFF;
            15'd3457: data <= 8'hFF;
            15'd3458: data <= 8'hFF;
            15'd3459: data <= 8'hFF;
            15'd3460: data <= 8'hFF;
            15'd3461: data <= 8'hFF;
            15'd3462: data <= 8'h00;
            15'd3463: data <= 8'h00;
            15'd3464: data <= 8'h3F;
            15'd3465: data <= 8'hFF;
            15'd3466: data <= 8'hC7;
            15'd3467: data <= 8'hFF;
            15'd3468: data <= 8'hFF;
            15'd3469: data <= 8'hFF;
            15'd3470: data <= 8'hFF;
            15'd3471: data <= 8'hFF;
            15'd3472: data <= 8'hFF;
            15'd3473: data <= 8'hFF;
            15'd3474: data <= 8'hFF;
            15'd3475: data <= 8'h80;
            15'd3476: data <= 8'h00;
            15'd3477: data <= 8'h00;
            15'd3478: data <= 8'h00;
            15'd3479: data <= 8'h00;
            15'd3480: data <= 8'h00;
            15'd3481: data <= 8'h00;
            15'd3482: data <= 8'h00;
            15'd3483: data <= 8'h00;
            15'd3484: data <= 8'h01;
            15'd3485: data <= 8'hFF;
            15'd3486: data <= 8'hFF;
            15'd3487: data <= 8'hFF;
            15'd3488: data <= 8'hFF;
            15'd3489: data <= 8'hFF;
            15'd3490: data <= 8'hFF;
            15'd3491: data <= 8'hFF;
            15'd3492: data <= 8'h00;
            15'd3493: data <= 8'h04;
            15'd3494: data <= 8'h3F;
            15'd3495: data <= 8'hFF;
            15'd3496: data <= 8'h8F;
            15'd3497: data <= 8'hFF;
            15'd3498: data <= 8'hFF;
            15'd3499: data <= 8'hFF;
            15'd3500: data <= 8'hFF;
            15'd3501: data <= 8'hFF;
            15'd3502: data <= 8'hFF;
            15'd3503: data <= 8'hFF;
            15'd3504: data <= 8'hFF;
            15'd3505: data <= 8'h80;
            15'd3506: data <= 8'h00;
            15'd3507: data <= 8'h00;
            15'd3508: data <= 8'h00;
            15'd3509: data <= 8'h00;
            15'd3510: data <= 8'h00;
            15'd3511: data <= 8'h00;
            15'd3512: data <= 8'h00;
            15'd3513: data <= 8'h00;
            15'd3514: data <= 8'h01;
            15'd3515: data <= 8'hFF;
            15'd3516: data <= 8'hFF;
            15'd3517: data <= 8'hFF;
            15'd3518: data <= 8'hFF;
            15'd3519: data <= 8'hFF;
            15'd3520: data <= 8'hFF;
            15'd3521: data <= 8'hFE;
            15'd3522: data <= 8'h0C;
            15'd3523: data <= 8'h1E;
            15'd3524: data <= 8'h3F;
            15'd3525: data <= 8'hFF;
            15'd3526: data <= 8'h9F;
            15'd3527: data <= 8'hFF;
            15'd3528: data <= 8'hFF;
            15'd3529: data <= 8'hFF;
            15'd3530: data <= 8'hFF;
            15'd3531: data <= 8'hFF;
            15'd3532: data <= 8'hFF;
            15'd3533: data <= 8'hFF;
            15'd3534: data <= 8'hFF;
            15'd3535: data <= 8'h80;
            15'd3536: data <= 8'h00;
            15'd3537: data <= 8'h00;
            15'd3538: data <= 8'h00;
            15'd3539: data <= 8'h00;
            15'd3540: data <= 8'h00;
            15'd3541: data <= 8'h00;
            15'd3542: data <= 8'h00;
            15'd3543: data <= 8'h00;
            15'd3544: data <= 8'h01;
            15'd3545: data <= 8'hFF;
            15'd3546: data <= 8'hFF;
            15'd3547: data <= 8'hFF;
            15'd3548: data <= 8'hFF;
            15'd3549: data <= 8'hFF;
            15'd3550: data <= 8'hFF;
            15'd3551: data <= 8'hFE;
            15'd3552: data <= 8'h1E;
            15'd3553: data <= 8'h3E;
            15'd3554: data <= 8'h3F;
            15'd3555: data <= 8'hFF;
            15'd3556: data <= 8'h3F;
            15'd3557: data <= 8'hFF;
            15'd3558: data <= 8'hFF;
            15'd3559: data <= 8'hFF;
            15'd3560: data <= 8'hFF;
            15'd3561: data <= 8'hFF;
            15'd3562: data <= 8'hFF;
            15'd3563: data <= 8'hFF;
            15'd3564: data <= 8'hFF;
            15'd3565: data <= 8'h80;
            15'd3566: data <= 8'h00;
            15'd3567: data <= 8'h00;
            15'd3568: data <= 8'h00;
            15'd3569: data <= 8'h00;
            15'd3570: data <= 8'h00;
            15'd3571: data <= 8'h00;
            15'd3572: data <= 8'h00;
            15'd3573: data <= 8'h00;
            15'd3574: data <= 8'h01;
            15'd3575: data <= 8'hFF;
            15'd3576: data <= 8'hFF;
            15'd3577: data <= 8'hFF;
            15'd3578: data <= 8'hFF;
            15'd3579: data <= 8'hFF;
            15'd3580: data <= 8'hFF;
            15'd3581: data <= 8'hFE;
            15'd3582: data <= 8'h1F;
            15'd3583: data <= 8'hFE;
            15'd3584: data <= 8'h3F;
            15'd3585: data <= 8'hFF;
            15'd3586: data <= 8'h3F;
            15'd3587: data <= 8'hFF;
            15'd3588: data <= 8'hFF;
            15'd3589: data <= 8'hFF;
            15'd3590: data <= 8'hFF;
            15'd3591: data <= 8'hFF;
            15'd3592: data <= 8'hFF;
            15'd3593: data <= 8'hFF;
            15'd3594: data <= 8'hFF;
            15'd3595: data <= 8'h80;
            15'd3596: data <= 8'h00;
            15'd3597: data <= 8'h00;
            15'd3598: data <= 8'h00;
            15'd3599: data <= 8'h00;
            15'd3600: data <= 8'h00;
            15'd3601: data <= 8'h00;
            15'd3602: data <= 8'h00;
            15'd3603: data <= 8'h00;
            15'd3604: data <= 8'h01;
            15'd3605: data <= 8'hFF;
            15'd3606: data <= 8'hFF;
            15'd3607: data <= 8'hFF;
            15'd3608: data <= 8'hFF;
            15'd3609: data <= 8'hFF;
            15'd3610: data <= 8'hFF;
            15'd3611: data <= 8'hFE;
            15'd3612: data <= 8'h1F;
            15'd3613: data <= 8'hFC;
            15'd3614: data <= 8'h3F;
            15'd3615: data <= 8'hFE;
            15'd3616: data <= 8'h7F;
            15'd3617: data <= 8'hFF;
            15'd3618: data <= 8'hFF;
            15'd3619: data <= 8'hFF;
            15'd3620: data <= 8'hFF;
            15'd3621: data <= 8'hFF;
            15'd3622: data <= 8'hFF;
            15'd3623: data <= 8'hFF;
            15'd3624: data <= 8'hFF;
            15'd3625: data <= 8'h80;
            15'd3626: data <= 8'h00;
            15'd3627: data <= 8'h00;
            15'd3628: data <= 8'h00;
            15'd3629: data <= 8'h00;
            15'd3630: data <= 8'h00;
            15'd3631: data <= 8'h00;
            15'd3632: data <= 8'h00;
            15'd3633: data <= 8'h00;
            15'd3634: data <= 8'h01;
            15'd3635: data <= 8'hFF;
            15'd3636: data <= 8'hFF;
            15'd3637: data <= 8'hFF;
            15'd3638: data <= 8'hFF;
            15'd3639: data <= 8'hFF;
            15'd3640: data <= 8'hFF;
            15'd3641: data <= 8'hFE;
            15'd3642: data <= 8'h1F;
            15'd3643: data <= 8'hFC;
            15'd3644: data <= 8'h3F;
            15'd3645: data <= 8'hFC;
            15'd3646: data <= 8'hFF;
            15'd3647: data <= 8'hFF;
            15'd3648: data <= 8'hFF;
            15'd3649: data <= 8'hFF;
            15'd3650: data <= 8'hFF;
            15'd3651: data <= 8'hFF;
            15'd3652: data <= 8'hFF;
            15'd3653: data <= 8'hFF;
            15'd3654: data <= 8'hFF;
            15'd3655: data <= 8'h80;
            15'd3656: data <= 8'h00;
            15'd3657: data <= 8'h00;
            15'd3658: data <= 8'h00;
            15'd3659: data <= 8'h00;
            15'd3660: data <= 8'h00;
            15'd3661: data <= 8'h00;
            15'd3662: data <= 8'h00;
            15'd3663: data <= 8'h00;
            15'd3664: data <= 8'h01;
            15'd3665: data <= 8'hFF;
            15'd3666: data <= 8'hFF;
            15'd3667: data <= 8'hFF;
            15'd3668: data <= 8'hFF;
            15'd3669: data <= 8'hFF;
            15'd3670: data <= 8'hFF;
            15'd3671: data <= 8'hFF;
            15'd3672: data <= 8'h0F;
            15'd3673: data <= 8'hF8;
            15'd3674: data <= 8'h7F;
            15'd3675: data <= 8'hFD;
            15'd3676: data <= 8'hFF;
            15'd3677: data <= 8'hFF;
            15'd3678: data <= 8'hFF;
            15'd3679: data <= 8'hFF;
            15'd3680: data <= 8'hFF;
            15'd3681: data <= 8'hFF;
            15'd3682: data <= 8'hFF;
            15'd3683: data <= 8'hFF;
            15'd3684: data <= 8'hFF;
            15'd3685: data <= 8'h80;
            15'd3686: data <= 8'h00;
            15'd3687: data <= 8'h00;
            15'd3688: data <= 8'h00;
            15'd3689: data <= 8'h00;
            15'd3690: data <= 8'h00;
            15'd3691: data <= 8'h00;
            15'd3692: data <= 8'h00;
            15'd3693: data <= 8'h00;
            15'd3694: data <= 8'h01;
            15'd3695: data <= 8'hFF;
            15'd3696: data <= 8'hFF;
            15'd3697: data <= 8'hFF;
            15'd3698: data <= 8'hFF;
            15'd3699: data <= 8'hFF;
            15'd3700: data <= 8'hFF;
            15'd3701: data <= 8'hFF;
            15'd3702: data <= 8'h87;
            15'd3703: data <= 8'hF8;
            15'd3704: data <= 8'h7F;
            15'd3705: data <= 8'hF9;
            15'd3706: data <= 8'hFF;
            15'd3707: data <= 8'hFF;
            15'd3708: data <= 8'hFF;
            15'd3709: data <= 8'hFF;
            15'd3710: data <= 8'hFF;
            15'd3711: data <= 8'hFF;
            15'd3712: data <= 8'hFF;
            15'd3713: data <= 8'hFF;
            15'd3714: data <= 8'hFF;
            15'd3715: data <= 8'h80;
            15'd3716: data <= 8'h00;
            15'd3717: data <= 8'h00;
            15'd3718: data <= 8'h00;
            15'd3719: data <= 8'h00;
            15'd3720: data <= 8'h00;
            15'd3721: data <= 8'h00;
            15'd3722: data <= 8'h00;
            15'd3723: data <= 8'h00;
            15'd3724: data <= 8'h01;
            15'd3725: data <= 8'hFF;
            15'd3726: data <= 8'hFF;
            15'd3727: data <= 8'hFF;
            15'd3728: data <= 8'hFF;
            15'd3729: data <= 8'hFF;
            15'd3730: data <= 8'hFF;
            15'd3731: data <= 8'hFF;
            15'd3732: data <= 8'h83;
            15'd3733: data <= 8'hF0;
            15'd3734: data <= 8'hFF;
            15'd3735: data <= 8'hFF;
            15'd3736: data <= 8'hFF;
            15'd3737: data <= 8'hFF;
            15'd3738: data <= 8'hFF;
            15'd3739: data <= 8'hFF;
            15'd3740: data <= 8'hFF;
            15'd3741: data <= 8'hFF;
            15'd3742: data <= 8'hFF;
            15'd3743: data <= 8'hFF;
            15'd3744: data <= 8'hFF;
            15'd3745: data <= 8'h80;
            15'd3746: data <= 8'h00;
            15'd3747: data <= 8'h00;
            15'd3748: data <= 8'h00;
            15'd3749: data <= 8'h00;
            15'd3750: data <= 8'h00;
            15'd3751: data <= 8'h00;
            15'd3752: data <= 8'h00;
            15'd3753: data <= 8'h00;
            15'd3754: data <= 8'h01;
            15'd3755: data <= 8'hFF;
            15'd3756: data <= 8'hFF;
            15'd3757: data <= 8'hFF;
            15'd3758: data <= 8'hFF;
            15'd3759: data <= 8'hFF;
            15'd3760: data <= 8'hFF;
            15'd3761: data <= 8'hFF;
            15'd3762: data <= 8'hC1;
            15'd3763: data <= 8'hE0;
            15'd3764: data <= 8'hFF;
            15'd3765: data <= 8'hFF;
            15'd3766: data <= 8'hFF;
            15'd3767: data <= 8'hFF;
            15'd3768: data <= 8'hFF;
            15'd3769: data <= 8'hFF;
            15'd3770: data <= 8'hFF;
            15'd3771: data <= 8'hFF;
            15'd3772: data <= 8'hFF;
            15'd3773: data <= 8'hFF;
            15'd3774: data <= 8'hFF;
            15'd3775: data <= 8'h80;
            15'd3776: data <= 8'h00;
            15'd3777: data <= 8'h00;
            15'd3778: data <= 8'h00;
            15'd3779: data <= 8'h00;
            15'd3780: data <= 8'h00;
            15'd3781: data <= 8'h00;
            15'd3782: data <= 8'h00;
            15'd3783: data <= 8'h00;
            15'd3784: data <= 8'h01;
            15'd3785: data <= 8'hFF;
            15'd3786: data <= 8'hFF;
            15'd3787: data <= 8'hFF;
            15'd3788: data <= 8'hFF;
            15'd3789: data <= 8'hFF;
            15'd3790: data <= 8'hFF;
            15'd3791: data <= 8'hFF;
            15'd3792: data <= 8'hE0;
            15'd3793: data <= 8'h41;
            15'd3794: data <= 8'hFF;
            15'd3795: data <= 8'hFF;
            15'd3796: data <= 8'hFF;
            15'd3797: data <= 8'hFF;
            15'd3798: data <= 8'hFF;
            15'd3799: data <= 8'hFF;
            15'd3800: data <= 8'hFF;
            15'd3801: data <= 8'hFF;
            15'd3802: data <= 8'hFF;
            15'd3803: data <= 8'hFF;
            15'd3804: data <= 8'hFF;
            15'd3805: data <= 8'h80;
            15'd3806: data <= 8'h00;
            15'd3807: data <= 8'h00;
            15'd3808: data <= 8'h00;
            15'd3809: data <= 8'h00;
            15'd3810: data <= 8'h00;
            15'd3811: data <= 8'h00;
            15'd3812: data <= 8'h00;
            15'd3813: data <= 8'h00;
            15'd3814: data <= 8'h01;
            15'd3815: data <= 8'hFF;
            15'd3816: data <= 8'hFF;
            15'd3817: data <= 8'hFF;
            15'd3818: data <= 8'hFF;
            15'd3819: data <= 8'hFF;
            15'd3820: data <= 8'hFF;
            15'd3821: data <= 8'hFF;
            15'd3822: data <= 8'hF8;
            15'd3823: data <= 8'h03;
            15'd3824: data <= 8'hFF;
            15'd3825: data <= 8'hFF;
            15'd3826: data <= 8'hFF;
            15'd3827: data <= 8'hFF;
            15'd3828: data <= 8'hFF;
            15'd3829: data <= 8'hFF;
            15'd3830: data <= 8'hFF;
            15'd3831: data <= 8'hFF;
            15'd3832: data <= 8'hFF;
            15'd3833: data <= 8'hFF;
            15'd3834: data <= 8'hFF;
            15'd3835: data <= 8'h80;
            15'd3836: data <= 8'h00;
            15'd3837: data <= 8'h00;
            15'd3838: data <= 8'h00;
            15'd3839: data <= 8'h00;
            15'd3840: data <= 8'h00;
            15'd3841: data <= 8'h00;
            15'd3842: data <= 8'h00;
            15'd3843: data <= 8'h00;
            15'd3844: data <= 8'h01;
            15'd3845: data <= 8'hFF;
            15'd3846: data <= 8'hFF;
            15'd3847: data <= 8'hFF;
            15'd3848: data <= 8'hFF;
            15'd3849: data <= 8'hFF;
            15'd3850: data <= 8'hFF;
            15'd3851: data <= 8'hFF;
            15'd3852: data <= 8'hEC;
            15'd3853: data <= 8'h07;
            15'd3854: data <= 8'hFF;
            15'd3855: data <= 8'hFF;
            15'd3856: data <= 8'hFF;
            15'd3857: data <= 8'hFF;
            15'd3858: data <= 8'hFF;
            15'd3859: data <= 8'hFF;
            15'd3860: data <= 8'hFF;
            15'd3861: data <= 8'hFF;
            15'd3862: data <= 8'hFF;
            15'd3863: data <= 8'hFF;
            15'd3864: data <= 8'hFF;
            15'd3865: data <= 8'h80;
            15'd3866: data <= 8'h00;
            15'd3867: data <= 8'h00;
            15'd3868: data <= 8'h00;
            15'd3869: data <= 8'h00;
            15'd3870: data <= 8'h00;
            15'd3871: data <= 8'h00;
            15'd3872: data <= 8'h00;
            15'd3873: data <= 8'h00;
            15'd3874: data <= 8'h01;
            15'd3875: data <= 8'hFF;
            15'd3876: data <= 8'hFF;
            15'd3877: data <= 8'hFF;
            15'd3878: data <= 8'hFF;
            15'd3879: data <= 8'hFF;
            15'd3880: data <= 8'hFF;
            15'd3881: data <= 8'hFF;
            15'd3882: data <= 8'hF6;
            15'd3883: data <= 8'h0F;
            15'd3884: data <= 8'hFF;
            15'd3885: data <= 8'hFF;
            15'd3886: data <= 8'hFF;
            15'd3887: data <= 8'hFF;
            15'd3888: data <= 8'hFF;
            15'd3889: data <= 8'hFF;
            15'd3890: data <= 8'hFF;
            15'd3891: data <= 8'hFF;
            15'd3892: data <= 8'hFF;
            15'd3893: data <= 8'hFF;
            15'd3894: data <= 8'hFF;
            15'd3895: data <= 8'h80;
            15'd3896: data <= 8'h00;
            15'd3897: data <= 8'h00;
            15'd3898: data <= 8'h00;
            15'd3899: data <= 8'h00;
            15'd3900: data <= 8'h00;
            15'd3901: data <= 8'h00;
            15'd3902: data <= 8'h00;
            15'd3903: data <= 8'h00;
            15'd3904: data <= 8'h01;
            15'd3905: data <= 8'hFF;
            15'd3906: data <= 8'hFD;
            15'd3907: data <= 8'hFF;
            15'd3908: data <= 8'hFF;
            15'd3909: data <= 8'hFF;
            15'd3910: data <= 8'hFF;
            15'd3911: data <= 8'hFF;
            15'd3912: data <= 8'hFF;
            15'd3913: data <= 8'hFF;
            15'd3914: data <= 8'hFF;
            15'd3915: data <= 8'hFF;
            15'd3916: data <= 8'hFF;
            15'd3917: data <= 8'hFF;
            15'd3918: data <= 8'hFF;
            15'd3919: data <= 8'hFF;
            15'd3920: data <= 8'hFF;
            15'd3921: data <= 8'hFF;
            15'd3922: data <= 8'hFF;
            15'd3923: data <= 8'hFF;
            15'd3924: data <= 8'hFF;
            15'd3925: data <= 8'h80;
            15'd3926: data <= 8'h00;
            15'd3927: data <= 8'h00;
            15'd3928: data <= 8'h00;
            15'd3929: data <= 8'h00;
            15'd3930: data <= 8'h00;
            15'd3931: data <= 8'h00;
            15'd3932: data <= 8'h00;
            15'd3933: data <= 8'h00;
            15'd3934: data <= 8'h01;
            15'd3935: data <= 8'hFF;
            15'd3936: data <= 8'hFF;
            15'd3937: data <= 8'hFF;
            15'd3938: data <= 8'hFF;
            15'd3939: data <= 8'hFF;
            15'd3940: data <= 8'hFF;
            15'd3941: data <= 8'hFF;
            15'd3942: data <= 8'hFF;
            15'd3943: data <= 8'hFF;
            15'd3944: data <= 8'hFF;
            15'd3945: data <= 8'hFF;
            15'd3946: data <= 8'hFF;
            15'd3947: data <= 8'hFF;
            15'd3948: data <= 8'hFF;
            15'd3949: data <= 8'hFF;
            15'd3950: data <= 8'hFF;
            15'd3951: data <= 8'hFF;
            15'd3952: data <= 8'hFF;
            15'd3953: data <= 8'hFF;
            15'd3954: data <= 8'hFF;
            15'd3955: data <= 8'h80;
            15'd3956: data <= 8'h00;
            15'd3957: data <= 8'h00;
            15'd3958: data <= 8'h00;
            15'd3959: data <= 8'h00;
            15'd3960: data <= 8'h00;
            15'd3961: data <= 8'h00;
            15'd3962: data <= 8'h00;
            15'd3963: data <= 8'h00;
            15'd3964: data <= 8'h01;
            15'd3965: data <= 8'hFF;
            15'd3966: data <= 8'hFF;
            15'd3967: data <= 8'hFF;
            15'd3968: data <= 8'hFF;
            15'd3969: data <= 8'hFF;
            15'd3970: data <= 8'hFF;
            15'd3971: data <= 8'hFF;
            15'd3972: data <= 8'hFF;
            15'd3973: data <= 8'hFF;
            15'd3974: data <= 8'hFF;
            15'd3975: data <= 8'hFF;
            15'd3976: data <= 8'hFF;
            15'd3977: data <= 8'hFF;
            15'd3978: data <= 8'hFF;
            15'd3979: data <= 8'hFF;
            15'd3980: data <= 8'hFF;
            15'd3981: data <= 8'hFF;
            15'd3982: data <= 8'hFF;
            15'd3983: data <= 8'hFF;
            15'd3984: data <= 8'hFF;
            15'd3985: data <= 8'h80;
            15'd3986: data <= 8'h00;
            15'd3987: data <= 8'h00;
            15'd3988: data <= 8'h00;
            15'd3989: data <= 8'h00;
            15'd3990: data <= 8'h00;
            15'd3991: data <= 8'h00;
            15'd3992: data <= 8'h00;
            15'd3993: data <= 8'h00;
            15'd3994: data <= 8'h01;
            15'd3995: data <= 8'hFF;
            15'd3996: data <= 8'hFF;
            15'd3997: data <= 8'hFF;
            15'd3998: data <= 8'hFF;
            15'd3999: data <= 8'hFF;
            15'd4000: data <= 8'hFF;
            15'd4001: data <= 8'hFF;
            15'd4002: data <= 8'hFF;
            15'd4003: data <= 8'hFF;
            15'd4004: data <= 8'hFF;
            15'd4005: data <= 8'hFF;
            15'd4006: data <= 8'hFF;
            15'd4007: data <= 8'hFF;
            15'd4008: data <= 8'hFF;
            15'd4009: data <= 8'hFF;
            15'd4010: data <= 8'hFF;
            15'd4011: data <= 8'hFF;
            15'd4012: data <= 8'hFF;
            15'd4013: data <= 8'hFF;
            15'd4014: data <= 8'hFF;
            15'd4015: data <= 8'h80;
            15'd4016: data <= 8'h00;
            15'd4017: data <= 8'h00;
            15'd4018: data <= 8'h00;
            15'd4019: data <= 8'h00;
            15'd4020: data <= 8'h00;
            15'd4021: data <= 8'h00;
            15'd4022: data <= 8'h00;
            15'd4023: data <= 8'h00;
            15'd4024: data <= 8'h01;
            15'd4025: data <= 8'hFF;
            15'd4026: data <= 8'hFF;
            15'd4027: data <= 8'hFF;
            15'd4028: data <= 8'hFF;
            15'd4029: data <= 8'hFF;
            15'd4030: data <= 8'hFF;
            15'd4031: data <= 8'hFF;
            15'd4032: data <= 8'hFF;
            15'd4033: data <= 8'hFF;
            15'd4034: data <= 8'hFF;
            15'd4035: data <= 8'hFF;
            15'd4036: data <= 8'hFF;
            15'd4037: data <= 8'hFF;
            15'd4038: data <= 8'hFF;
            15'd4039: data <= 8'hFF;
            15'd4040: data <= 8'hFF;
            15'd4041: data <= 8'hFF;
            15'd4042: data <= 8'hFF;
            15'd4043: data <= 8'hFF;
            15'd4044: data <= 8'hFF;
            15'd4045: data <= 8'h80;
            15'd4046: data <= 8'h00;
            15'd4047: data <= 8'h00;
            15'd4048: data <= 8'h00;
            15'd4049: data <= 8'h00;
            15'd4050: data <= 8'h00;
            15'd4051: data <= 8'h00;
            15'd4052: data <= 8'h00;
            15'd4053: data <= 8'h00;
            15'd4054: data <= 8'h01;
            15'd4055: data <= 8'hFF;
            15'd4056: data <= 8'hFF;
            15'd4057: data <= 8'hFF;
            15'd4058: data <= 8'hFF;
            15'd4059: data <= 8'hFF;
            15'd4060: data <= 8'hFF;
            15'd4061: data <= 8'hFF;
            15'd4062: data <= 8'hFF;
            15'd4063: data <= 8'hFF;
            15'd4064: data <= 8'hFF;
            15'd4065: data <= 8'hFF;
            15'd4066: data <= 8'hFF;
            15'd4067: data <= 8'hFF;
            15'd4068: data <= 8'hFF;
            15'd4069: data <= 8'hFF;
            15'd4070: data <= 8'hFF;
            15'd4071: data <= 8'hFF;
            15'd4072: data <= 8'hFF;
            15'd4073: data <= 8'hFF;
            15'd4074: data <= 8'hFF;
            15'd4075: data <= 8'h80;
            15'd4076: data <= 8'h00;
            15'd4077: data <= 8'h00;
            15'd4078: data <= 8'h00;
            15'd4079: data <= 8'h00;
            15'd4080: data <= 8'h00;
            15'd4081: data <= 8'h00;
            15'd4082: data <= 8'h00;
            15'd4083: data <= 8'h00;
            15'd4084: data <= 8'h01;
            15'd4085: data <= 8'hFF;
            15'd4086: data <= 8'hFF;
            15'd4087: data <= 8'hFF;
            15'd4088: data <= 8'hFF;
            15'd4089: data <= 8'hFF;
            15'd4090: data <= 8'hFF;
            15'd4091: data <= 8'hFF;
            15'd4092: data <= 8'hFF;
            15'd4093: data <= 8'hFF;
            15'd4094: data <= 8'hFF;
            15'd4095: data <= 8'hFF;
            15'd4096: data <= 8'hFF;
            15'd4097: data <= 8'hFF;
            15'd4098: data <= 8'hFF;
            15'd4099: data <= 8'hFF;
            15'd4100: data <= 8'hFF;
            15'd4101: data <= 8'hFF;
            15'd4102: data <= 8'hFF;
            15'd4103: data <= 8'hFF;
            15'd4104: data <= 8'hFF;
            15'd4105: data <= 8'h80;
            15'd4106: data <= 8'h00;
            15'd4107: data <= 8'h00;
            15'd4108: data <= 8'h00;
            15'd4109: data <= 8'h00;
            15'd4110: data <= 8'h00;
            15'd4111: data <= 8'h00;
            15'd4112: data <= 8'h00;
            15'd4113: data <= 8'h00;
            15'd4114: data <= 8'h01;
            15'd4115: data <= 8'hFF;
            15'd4116: data <= 8'hFF;
            15'd4117: data <= 8'hFF;
            15'd4118: data <= 8'hFF;
            15'd4119: data <= 8'hFF;
            15'd4120: data <= 8'hFF;
            15'd4121: data <= 8'hFF;
            15'd4122: data <= 8'hFF;
            15'd4123: data <= 8'hFF;
            15'd4124: data <= 8'hFF;
            15'd4125: data <= 8'hFF;
            15'd4126: data <= 8'hFF;
            15'd4127: data <= 8'hFF;
            15'd4128: data <= 8'hFF;
            15'd4129: data <= 8'hFF;
            15'd4130: data <= 8'hFF;
            15'd4131: data <= 8'hFF;
            15'd4132: data <= 8'hFF;
            15'd4133: data <= 8'hFF;
            15'd4134: data <= 8'hFF;
            15'd4135: data <= 8'h80;
            15'd4136: data <= 8'h00;
            15'd4137: data <= 8'h00;
            15'd4138: data <= 8'h00;
            15'd4139: data <= 8'h00;
            15'd4140: data <= 8'h00;
            15'd4141: data <= 8'h00;
            15'd4142: data <= 8'h00;
            15'd4143: data <= 8'h00;
            15'd4144: data <= 8'h01;
            15'd4145: data <= 8'hFF;
            15'd4146: data <= 8'hFF;
            15'd4147: data <= 8'hFF;
            15'd4148: data <= 8'hFF;
            15'd4149: data <= 8'hFF;
            15'd4150: data <= 8'hFF;
            15'd4151: data <= 8'hFF;
            15'd4152: data <= 8'hFF;
            15'd4153: data <= 8'hFF;
            15'd4154: data <= 8'hFF;
            15'd4155: data <= 8'hFF;
            15'd4156: data <= 8'hFF;
            15'd4157: data <= 8'hFF;
            15'd4158: data <= 8'hFF;
            15'd4159: data <= 8'hFF;
            15'd4160: data <= 8'hFF;
            15'd4161: data <= 8'hFF;
            15'd4162: data <= 8'hFF;
            15'd4163: data <= 8'hFF;
            15'd4164: data <= 8'hFF;
            15'd4165: data <= 8'h80;
            15'd4166: data <= 8'h00;
            15'd4167: data <= 8'h00;
            15'd4168: data <= 8'h00;
            15'd4169: data <= 8'h00;
            15'd4170: data <= 8'h00;
            15'd4171: data <= 8'h00;
            15'd4172: data <= 8'h00;
            15'd4173: data <= 8'h00;
            15'd4174: data <= 8'h01;
            15'd4175: data <= 8'hFF;
            15'd4176: data <= 8'hFF;
            15'd4177: data <= 8'hFF;
            15'd4178: data <= 8'hFF;
            15'd4179: data <= 8'hFF;
            15'd4180: data <= 8'hFF;
            15'd4181: data <= 8'hFF;
            15'd4182: data <= 8'hFF;
            15'd4183: data <= 8'hFF;
            15'd4184: data <= 8'hFF;
            15'd4185: data <= 8'hFF;
            15'd4186: data <= 8'hFF;
            15'd4187: data <= 8'hFF;
            15'd4188: data <= 8'hFF;
            15'd4189: data <= 8'hFF;
            15'd4190: data <= 8'hFF;
            15'd4191: data <= 8'hFF;
            15'd4192: data <= 8'hFF;
            15'd4193: data <= 8'hFF;
            15'd4194: data <= 8'hFF;
            15'd4195: data <= 8'h80;
            15'd4196: data <= 8'h00;
            15'd4197: data <= 8'h00;
            15'd4198: data <= 8'h00;
            15'd4199: data <= 8'h00;
            15'd4200: data <= 8'h00;
            15'd4201: data <= 8'h00;
            15'd4202: data <= 8'h00;
            15'd4203: data <= 8'h00;
            15'd4204: data <= 8'h01;
            15'd4205: data <= 8'hFF;
            15'd4206: data <= 8'hFF;
            15'd4207: data <= 8'hFF;
            15'd4208: data <= 8'hFF;
            15'd4209: data <= 8'hFF;
            15'd4210: data <= 8'hFF;
            15'd4211: data <= 8'hFF;
            15'd4212: data <= 8'hFF;
            15'd4213: data <= 8'hFF;
            15'd4214: data <= 8'hFF;
            15'd4215: data <= 8'hFF;
            15'd4216: data <= 8'hFF;
            15'd4217: data <= 8'hFF;
            15'd4218: data <= 8'hFF;
            15'd4219: data <= 8'hFF;
            15'd4220: data <= 8'hFF;
            15'd4221: data <= 8'hFF;
            15'd4222: data <= 8'hFF;
            15'd4223: data <= 8'hFF;
            15'd4224: data <= 8'hFF;
            15'd4225: data <= 8'h80;
            15'd4226: data <= 8'h00;
            15'd4227: data <= 8'h00;
            15'd4228: data <= 8'h00;
            15'd4229: data <= 8'h00;
            15'd4230: data <= 8'h00;
            15'd4231: data <= 8'h00;
            15'd4232: data <= 8'h00;
            15'd4233: data <= 8'h00;
            15'd4234: data <= 8'h01;
            15'd4235: data <= 8'hFF;
            15'd4236: data <= 8'hFF;
            15'd4237: data <= 8'hFF;
            15'd4238: data <= 8'hFF;
            15'd4239: data <= 8'hFF;
            15'd4240: data <= 8'hFF;
            15'd4241: data <= 8'hFF;
            15'd4242: data <= 8'hFF;
            15'd4243: data <= 8'hFF;
            15'd4244: data <= 8'hFF;
            15'd4245: data <= 8'hFF;
            15'd4246: data <= 8'hFF;
            15'd4247: data <= 8'hFF;
            15'd4248: data <= 8'hFF;
            15'd4249: data <= 8'hFF;
            15'd4250: data <= 8'hFF;
            15'd4251: data <= 8'hFF;
            15'd4252: data <= 8'hFF;
            15'd4253: data <= 8'hFF;
            15'd4254: data <= 8'hFF;
            15'd4255: data <= 8'h80;
            15'd4256: data <= 8'h00;
            15'd4257: data <= 8'h00;
            15'd4258: data <= 8'h00;
            15'd4259: data <= 8'h00;
            15'd4260: data <= 8'h00;
            15'd4261: data <= 8'h00;
            15'd4262: data <= 8'h00;
            15'd4263: data <= 8'h00;
            15'd4264: data <= 8'h01;
            15'd4265: data <= 8'hFF;
            15'd4266: data <= 8'hFF;
            15'd4267: data <= 8'hFF;
            15'd4268: data <= 8'hFF;
            15'd4269: data <= 8'hFF;
            15'd4270: data <= 8'hFF;
            15'd4271: data <= 8'hFF;
            15'd4272: data <= 8'hFF;
            15'd4273: data <= 8'hFF;
            15'd4274: data <= 8'hFF;
            15'd4275: data <= 8'hFF;
            15'd4276: data <= 8'hFF;
            15'd4277: data <= 8'hFF;
            15'd4278: data <= 8'hFF;
            15'd4279: data <= 8'hFF;
            15'd4280: data <= 8'hFF;
            15'd4281: data <= 8'hFF;
            15'd4282: data <= 8'hFF;
            15'd4283: data <= 8'hFF;
            15'd4284: data <= 8'hFF;
            15'd4285: data <= 8'h80;
            15'd4286: data <= 8'h00;
            15'd4287: data <= 8'h00;
            15'd4288: data <= 8'h00;
            15'd4289: data <= 8'h00;
            15'd4290: data <= 8'h00;
            15'd4291: data <= 8'h00;
            15'd4292: data <= 8'h00;
            15'd4293: data <= 8'h00;
            15'd4294: data <= 8'h01;
            15'd4295: data <= 8'hFF;
            15'd4296: data <= 8'hFF;
            15'd4297: data <= 8'hFF;
            15'd4298: data <= 8'hFF;
            15'd4299: data <= 8'hFF;
            15'd4300: data <= 8'hFF;
            15'd4301: data <= 8'hFF;
            15'd4302: data <= 8'hFF;
            15'd4303: data <= 8'hFF;
            15'd4304: data <= 8'hFF;
            15'd4305: data <= 8'hFF;
            15'd4306: data <= 8'hFF;
            15'd4307: data <= 8'hFF;
            15'd4308: data <= 8'hFF;
            15'd4309: data <= 8'hFF;
            15'd4310: data <= 8'hFF;
            15'd4311: data <= 8'hFF;
            15'd4312: data <= 8'hFF;
            15'd4313: data <= 8'hFF;
            15'd4314: data <= 8'hFF;
            15'd4315: data <= 8'h80;
            15'd4316: data <= 8'h00;
            15'd4317: data <= 8'h00;
            15'd4318: data <= 8'h00;
            15'd4319: data <= 8'h00;
            15'd4320: data <= 8'h00;
            15'd4321: data <= 8'h00;
            15'd4322: data <= 8'h00;
            15'd4323: data <= 8'h00;
            15'd4324: data <= 8'h01;
            15'd4325: data <= 8'hFF;
            15'd4326: data <= 8'hFF;
            15'd4327: data <= 8'hFF;
            15'd4328: data <= 8'hFF;
            15'd4329: data <= 8'hFF;
            15'd4330: data <= 8'hFF;
            15'd4331: data <= 8'hFF;
            15'd4332: data <= 8'hFF;
            15'd4333: data <= 8'hEF;
            15'd4334: data <= 8'hFF;
            15'd4335: data <= 8'hF3;
            15'd4336: data <= 8'hFF;
            15'd4337: data <= 8'hFF;
            15'd4338: data <= 8'hFF;
            15'd4339: data <= 8'hFF;
            15'd4340: data <= 8'hFF;
            15'd4341: data <= 8'hFF;
            15'd4342: data <= 8'hFF;
            15'd4343: data <= 8'hFF;
            15'd4344: data <= 8'hFF;
            15'd4345: data <= 8'h80;
            15'd4346: data <= 8'h00;
            15'd4347: data <= 8'h00;
            15'd4348: data <= 8'h00;
            15'd4349: data <= 8'h00;
            15'd4350: data <= 8'h00;
            15'd4351: data <= 8'h00;
            15'd4352: data <= 8'h00;
            15'd4353: data <= 8'h00;
            15'd4354: data <= 8'h01;
            15'd4355: data <= 8'hFF;
            15'd4356: data <= 8'hFF;
            15'd4357: data <= 8'hFF;
            15'd4358: data <= 8'hFF;
            15'd4359: data <= 8'hFF;
            15'd4360: data <= 8'hFF;
            15'd4361: data <= 8'hFF;
            15'd4362: data <= 8'hFC;
            15'd4363: data <= 8'hC7;
            15'd4364: data <= 8'hFF;
            15'd4365: data <= 8'hF0;
            15'd4366: data <= 8'h03;
            15'd4367: data <= 8'hFF;
            15'd4368: data <= 8'hFF;
            15'd4369: data <= 8'hFF;
            15'd4370: data <= 8'hFF;
            15'd4371: data <= 8'hFF;
            15'd4372: data <= 8'hFF;
            15'd4373: data <= 8'hFF;
            15'd4374: data <= 8'hFF;
            15'd4375: data <= 8'h80;
            15'd4376: data <= 8'h00;
            15'd4377: data <= 8'h00;
            15'd4378: data <= 8'h00;
            15'd4379: data <= 8'h00;
            15'd4380: data <= 8'h00;
            15'd4381: data <= 8'h00;
            15'd4382: data <= 8'h00;
            15'd4383: data <= 8'h00;
            15'd4384: data <= 8'h01;
            15'd4385: data <= 8'hFF;
            15'd4386: data <= 8'hFF;
            15'd4387: data <= 8'hFF;
            15'd4388: data <= 8'hFF;
            15'd4389: data <= 8'hFF;
            15'd4390: data <= 8'hFF;
            15'd4391: data <= 8'hFF;
            15'd4392: data <= 8'hFC;
            15'd4393: data <= 8'h47;
            15'd4394: data <= 8'hFF;
            15'd4395: data <= 8'hE0;
            15'd4396: data <= 8'h01;
            15'd4397: data <= 8'hFF;
            15'd4398: data <= 8'hFF;
            15'd4399: data <= 8'hFF;
            15'd4400: data <= 8'hFF;
            15'd4401: data <= 8'hFF;
            15'd4402: data <= 8'hFF;
            15'd4403: data <= 8'hFF;
            15'd4404: data <= 8'hFF;
            15'd4405: data <= 8'h80;
            15'd4406: data <= 8'h00;
            15'd4407: data <= 8'h00;
            15'd4408: data <= 8'h00;
            15'd4409: data <= 8'h00;
            15'd4410: data <= 8'h00;
            15'd4411: data <= 8'h00;
            15'd4412: data <= 8'h00;
            15'd4413: data <= 8'h00;
            15'd4414: data <= 8'h01;
            15'd4415: data <= 8'hFF;
            15'd4416: data <= 8'hFF;
            15'd4417: data <= 8'hFF;
            15'd4418: data <= 8'hFF;
            15'd4419: data <= 8'hFF;
            15'd4420: data <= 8'hFF;
            15'd4421: data <= 8'hFF;
            15'd4422: data <= 8'hFC;
            15'd4423: data <= 8'hC0;
            15'd4424: data <= 8'h7F;
            15'd4425: data <= 8'hE0;
            15'd4426: data <= 8'h03;
            15'd4427: data <= 8'hFF;
            15'd4428: data <= 8'hF3;
            15'd4429: data <= 8'hFF;
            15'd4430: data <= 8'hFF;
            15'd4431: data <= 8'hFF;
            15'd4432: data <= 8'hFF;
            15'd4433: data <= 8'hFF;
            15'd4434: data <= 8'hFF;
            15'd4435: data <= 8'h80;
            15'd4436: data <= 8'h00;
            15'd4437: data <= 8'h00;
            15'd4438: data <= 8'h00;
            15'd4439: data <= 8'h00;
            15'd4440: data <= 8'h00;
            15'd4441: data <= 8'h00;
            15'd4442: data <= 8'h00;
            15'd4443: data <= 8'h00;
            15'd4444: data <= 8'h01;
            15'd4445: data <= 8'hFF;
            15'd4446: data <= 8'hFF;
            15'd4447: data <= 8'hFF;
            15'd4448: data <= 8'hFF;
            15'd4449: data <= 8'hFF;
            15'd4450: data <= 8'hFF;
            15'd4451: data <= 8'hFF;
            15'd4452: data <= 8'hF8;
            15'd4453: data <= 8'h00;
            15'd4454: data <= 8'h7F;
            15'd4455: data <= 8'hC7;
            15'd4456: data <= 8'hFF;
            15'd4457: data <= 8'hFF;
            15'd4458: data <= 8'hF1;
            15'd4459: data <= 8'hFF;
            15'd4460: data <= 8'hFF;
            15'd4461: data <= 8'hFF;
            15'd4462: data <= 8'hFF;
            15'd4463: data <= 8'hFF;
            15'd4464: data <= 8'hFF;
            15'd4465: data <= 8'h80;
            15'd4466: data <= 8'h00;
            15'd4467: data <= 8'h00;
            15'd4468: data <= 8'h00;
            15'd4469: data <= 8'h00;
            15'd4470: data <= 8'h00;
            15'd4471: data <= 8'h00;
            15'd4472: data <= 8'h00;
            15'd4473: data <= 8'h00;
            15'd4474: data <= 8'h01;
            15'd4475: data <= 8'hFF;
            15'd4476: data <= 8'hFF;
            15'd4477: data <= 8'hFF;
            15'd4478: data <= 8'hFF;
            15'd4479: data <= 8'hFF;
            15'd4480: data <= 8'hFF;
            15'd4481: data <= 8'hFF;
            15'd4482: data <= 8'hF8;
            15'd4483: data <= 8'h00;
            15'd4484: data <= 8'hFF;
            15'd4485: data <= 8'h80;
            15'd4486: data <= 8'h03;
            15'd4487: data <= 8'hFF;
            15'd4488: data <= 8'hE1;
            15'd4489: data <= 8'hFF;
            15'd4490: data <= 8'hFF;
            15'd4491: data <= 8'hFF;
            15'd4492: data <= 8'hFF;
            15'd4493: data <= 8'hFF;
            15'd4494: data <= 8'hFF;
            15'd4495: data <= 8'h80;
            15'd4496: data <= 8'h00;
            15'd4497: data <= 8'h00;
            15'd4498: data <= 8'h00;
            15'd4499: data <= 8'h00;
            15'd4500: data <= 8'h00;
            15'd4501: data <= 8'h00;
            15'd4502: data <= 8'h00;
            15'd4503: data <= 8'h00;
            15'd4504: data <= 8'h01;
            15'd4505: data <= 8'hFF;
            15'd4506: data <= 8'hFF;
            15'd4507: data <= 8'hFF;
            15'd4508: data <= 8'hFF;
            15'd4509: data <= 8'hFF;
            15'd4510: data <= 8'hFF;
            15'd4511: data <= 8'hFF;
            15'd4512: data <= 8'hF8;
            15'd4513: data <= 8'hC7;
            15'd4514: data <= 8'hFF;
            15'd4515: data <= 8'h88;
            15'd4516: data <= 8'h03;
            15'd4517: data <= 8'hFF;
            15'd4518: data <= 8'hE3;
            15'd4519: data <= 8'hFF;
            15'd4520: data <= 8'hFF;
            15'd4521: data <= 8'hFF;
            15'd4522: data <= 8'hFF;
            15'd4523: data <= 8'hFF;
            15'd4524: data <= 8'hFF;
            15'd4525: data <= 8'h80;
            15'd4526: data <= 8'h00;
            15'd4527: data <= 8'h00;
            15'd4528: data <= 8'h00;
            15'd4529: data <= 8'h00;
            15'd4530: data <= 8'h00;
            15'd4531: data <= 8'h00;
            15'd4532: data <= 8'h00;
            15'd4533: data <= 8'h00;
            15'd4534: data <= 8'h01;
            15'd4535: data <= 8'hFF;
            15'd4536: data <= 8'hFF;
            15'd4537: data <= 8'hFF;
            15'd4538: data <= 8'hFF;
            15'd4539: data <= 8'hFF;
            15'd4540: data <= 8'hFF;
            15'd4541: data <= 8'hFF;
            15'd4542: data <= 8'hF1;
            15'd4543: data <= 8'h87;
            15'd4544: data <= 8'hFF;
            15'd4545: data <= 8'h9F;
            15'd4546: data <= 8'hFF;
            15'd4547: data <= 8'hFF;
            15'd4548: data <= 8'hE3;
            15'd4549: data <= 8'hFF;
            15'd4550: data <= 8'hFF;
            15'd4551: data <= 8'hFF;
            15'd4552: data <= 8'hFF;
            15'd4553: data <= 8'hFF;
            15'd4554: data <= 8'hFF;
            15'd4555: data <= 8'h80;
            15'd4556: data <= 8'h00;
            15'd4557: data <= 8'h00;
            15'd4558: data <= 8'h00;
            15'd4559: data <= 8'h00;
            15'd4560: data <= 8'h00;
            15'd4561: data <= 8'h00;
            15'd4562: data <= 8'h00;
            15'd4563: data <= 8'h00;
            15'd4564: data <= 8'h01;
            15'd4565: data <= 8'hFF;
            15'd4566: data <= 8'hFF;
            15'd4567: data <= 8'hFF;
            15'd4568: data <= 8'hFF;
            15'd4569: data <= 8'hFF;
            15'd4570: data <= 8'hFF;
            15'd4571: data <= 8'hFF;
            15'd4572: data <= 8'hF1;
            15'd4573: data <= 8'hC7;
            15'd4574: data <= 8'hFF;
            15'd4575: data <= 8'hF8;
            15'd4576: data <= 8'h01;
            15'd4577: data <= 8'hFF;
            15'd4578: data <= 8'hE3;
            15'd4579: data <= 8'hFF;
            15'd4580: data <= 8'hFF;
            15'd4581: data <= 8'hFF;
            15'd4582: data <= 8'hFF;
            15'd4583: data <= 8'hFF;
            15'd4584: data <= 8'hFF;
            15'd4585: data <= 8'h80;
            15'd4586: data <= 8'h00;
            15'd4587: data <= 8'h00;
            15'd4588: data <= 8'h00;
            15'd4589: data <= 8'h00;
            15'd4590: data <= 8'h00;
            15'd4591: data <= 8'h00;
            15'd4592: data <= 8'h00;
            15'd4593: data <= 8'h00;
            15'd4594: data <= 8'h01;
            15'd4595: data <= 8'hFF;
            15'd4596: data <= 8'hFF;
            15'd4597: data <= 8'hFF;
            15'd4598: data <= 8'hFF;
            15'd4599: data <= 8'hFF;
            15'd4600: data <= 8'hFF;
            15'd4601: data <= 8'hFF;
            15'd4602: data <= 8'hF3;
            15'd4603: data <= 8'hC1;
            15'd4604: data <= 8'hFF;
            15'd4605: data <= 8'hF0;
            15'd4606: data <= 8'h01;
            15'd4607: data <= 8'hFF;
            15'd4608: data <= 8'hF3;
            15'd4609: data <= 8'hFF;
            15'd4610: data <= 8'hFF;
            15'd4611: data <= 8'hFF;
            15'd4612: data <= 8'hFF;
            15'd4613: data <= 8'hFF;
            15'd4614: data <= 8'hFF;
            15'd4615: data <= 8'h80;
            15'd4616: data <= 8'h00;
            15'd4617: data <= 8'h00;
            15'd4618: data <= 8'h00;
            15'd4619: data <= 8'h00;
            15'd4620: data <= 8'h00;
            15'd4621: data <= 8'h00;
            15'd4622: data <= 8'h00;
            15'd4623: data <= 8'h00;
            15'd4624: data <= 8'h01;
            15'd4625: data <= 8'hFF;
            15'd4626: data <= 8'hFF;
            15'd4627: data <= 8'hFF;
            15'd4628: data <= 8'hFF;
            15'd4629: data <= 8'hFF;
            15'd4630: data <= 8'hFF;
            15'd4631: data <= 8'hFF;
            15'd4632: data <= 8'hFE;
            15'd4633: data <= 8'h00;
            15'd4634: data <= 8'h7F;
            15'd4635: data <= 8'hF8;
            15'd4636: data <= 8'h11;
            15'd4637: data <= 8'hFF;
            15'd4638: data <= 8'hF3;
            15'd4639: data <= 8'hFF;
            15'd4640: data <= 8'hFF;
            15'd4641: data <= 8'hFF;
            15'd4642: data <= 8'hFF;
            15'd4643: data <= 8'hFF;
            15'd4644: data <= 8'hFF;
            15'd4645: data <= 8'h80;
            15'd4646: data <= 8'h00;
            15'd4647: data <= 8'h00;
            15'd4648: data <= 8'h00;
            15'd4649: data <= 8'h00;
            15'd4650: data <= 8'h00;
            15'd4651: data <= 8'h00;
            15'd4652: data <= 8'h00;
            15'd4653: data <= 8'h00;
            15'd4654: data <= 8'h01;
            15'd4655: data <= 8'hFF;
            15'd4656: data <= 8'hFF;
            15'd4657: data <= 8'hFF;
            15'd4658: data <= 8'hFF;
            15'd4659: data <= 8'hFF;
            15'd4660: data <= 8'hFF;
            15'd4661: data <= 8'hFF;
            15'd4662: data <= 8'hFC;
            15'd4663: data <= 8'h00;
            15'd4664: data <= 8'h7F;
            15'd4665: data <= 8'hFF;
            15'd4666: data <= 8'hF9;
            15'd4667: data <= 8'hFF;
            15'd4668: data <= 8'hF3;
            15'd4669: data <= 8'hFF;
            15'd4670: data <= 8'hFF;
            15'd4671: data <= 8'hFF;
            15'd4672: data <= 8'hFF;
            15'd4673: data <= 8'hFF;
            15'd4674: data <= 8'hFF;
            15'd4675: data <= 8'h80;
            15'd4676: data <= 8'h00;
            15'd4677: data <= 8'h00;
            15'd4678: data <= 8'h00;
            15'd4679: data <= 8'h00;
            15'd4680: data <= 8'h00;
            15'd4681: data <= 8'h00;
            15'd4682: data <= 8'h00;
            15'd4683: data <= 8'h00;
            15'd4684: data <= 8'h01;
            15'd4685: data <= 8'hFF;
            15'd4686: data <= 8'hFF;
            15'd4687: data <= 8'hFF;
            15'd4688: data <= 8'hFF;
            15'd4689: data <= 8'hFF;
            15'd4690: data <= 8'hFF;
            15'd4691: data <= 8'hFF;
            15'd4692: data <= 8'hFE;
            15'd4693: data <= 8'h03;
            15'd4694: data <= 8'hFF;
            15'd4695: data <= 8'hFF;
            15'd4696: data <= 8'hF9;
            15'd4697: data <= 8'hFF;
            15'd4698: data <= 8'hFF;
            15'd4699: data <= 8'hFF;
            15'd4700: data <= 8'hFF;
            15'd4701: data <= 8'hFF;
            15'd4702: data <= 8'hFF;
            15'd4703: data <= 8'hFF;
            15'd4704: data <= 8'hFF;
            15'd4705: data <= 8'h80;
            15'd4706: data <= 8'h00;
            15'd4707: data <= 8'h00;
            15'd4708: data <= 8'h00;
            15'd4709: data <= 8'h00;
            15'd4710: data <= 8'h00;
            15'd4711: data <= 8'h00;
            15'd4712: data <= 8'h00;
            15'd4713: data <= 8'h00;
            15'd4714: data <= 8'h01;
            15'd4715: data <= 8'hFF;
            15'd4716: data <= 8'hFF;
            15'd4717: data <= 8'hFF;
            15'd4718: data <= 8'hFF;
            15'd4719: data <= 8'hFF;
            15'd4720: data <= 8'hFF;
            15'd4721: data <= 8'hFF;
            15'd4722: data <= 8'hFF;
            15'd4723: data <= 8'hC7;
            15'd4724: data <= 8'hFF;
            15'd4725: data <= 8'hFF;
            15'd4726: data <= 8'hF8;
            15'd4727: data <= 8'hFF;
            15'd4728: data <= 8'hFF;
            15'd4729: data <= 8'hFF;
            15'd4730: data <= 8'hFF;
            15'd4731: data <= 8'hFF;
            15'd4732: data <= 8'hFF;
            15'd4733: data <= 8'hFF;
            15'd4734: data <= 8'hFF;
            15'd4735: data <= 8'h80;
            15'd4736: data <= 8'h00;
            15'd4737: data <= 8'h00;
            15'd4738: data <= 8'h00;
            15'd4739: data <= 8'h00;
            15'd4740: data <= 8'h00;
            15'd4741: data <= 8'h00;
            15'd4742: data <= 8'h00;
            15'd4743: data <= 8'h00;
            15'd4744: data <= 8'h01;
            15'd4745: data <= 8'hFF;
            15'd4746: data <= 8'hFF;
            15'd4747: data <= 8'hFF;
            15'd4748: data <= 8'hFF;
            15'd4749: data <= 8'hFF;
            15'd4750: data <= 8'hFF;
            15'd4751: data <= 8'hFF;
            15'd4752: data <= 8'hFF;
            15'd4753: data <= 8'hC7;
            15'd4754: data <= 8'hFF;
            15'd4755: data <= 8'hFF;
            15'd4756: data <= 8'hF8;
            15'd4757: data <= 8'hBF;
            15'd4758: data <= 8'hE7;
            15'd4759: data <= 8'hFF;
            15'd4760: data <= 8'hFF;
            15'd4761: data <= 8'hFF;
            15'd4762: data <= 8'hFF;
            15'd4763: data <= 8'hFF;
            15'd4764: data <= 8'hFF;
            15'd4765: data <= 8'h80;
            15'd4766: data <= 8'h00;
            15'd4767: data <= 8'h00;
            15'd4768: data <= 8'h00;
            15'd4769: data <= 8'h00;
            15'd4770: data <= 8'h00;
            15'd4771: data <= 8'h00;
            15'd4772: data <= 8'h00;
            15'd4773: data <= 8'h00;
            15'd4774: data <= 8'h01;
            15'd4775: data <= 8'hFF;
            15'd4776: data <= 8'hFF;
            15'd4777: data <= 8'hFF;
            15'd4778: data <= 8'hFF;
            15'd4779: data <= 8'hFF;
            15'd4780: data <= 8'hFF;
            15'd4781: data <= 8'hFF;
            15'd4782: data <= 8'hF1;
            15'd4783: data <= 8'h00;
            15'd4784: data <= 8'h1F;
            15'd4785: data <= 8'hFF;
            15'd4786: data <= 8'hFC;
            15'd4787: data <= 8'h1F;
            15'd4788: data <= 8'hE3;
            15'd4789: data <= 8'hFF;
            15'd4790: data <= 8'hFF;
            15'd4791: data <= 8'hFF;
            15'd4792: data <= 8'hFF;
            15'd4793: data <= 8'hFF;
            15'd4794: data <= 8'hFF;
            15'd4795: data <= 8'h80;
            15'd4796: data <= 8'h00;
            15'd4797: data <= 8'h00;
            15'd4798: data <= 8'h00;
            15'd4799: data <= 8'h00;
            15'd4800: data <= 8'h00;
            15'd4801: data <= 8'h00;
            15'd4802: data <= 8'h00;
            15'd4803: data <= 8'h00;
            15'd4804: data <= 8'h01;
            15'd4805: data <= 8'hFF;
            15'd4806: data <= 8'hFF;
            15'd4807: data <= 8'hFF;
            15'd4808: data <= 8'hFF;
            15'd4809: data <= 8'hFF;
            15'd4810: data <= 8'hFF;
            15'd4811: data <= 8'hFF;
            15'd4812: data <= 8'hE0;
            15'd4813: data <= 8'h00;
            15'd4814: data <= 8'h0F;
            15'd4815: data <= 8'hFF;
            15'd4816: data <= 8'hFC;
            15'd4817: data <= 8'h1F;
            15'd4818: data <= 8'hE7;
            15'd4819: data <= 8'hFF;
            15'd4820: data <= 8'hFF;
            15'd4821: data <= 8'hFF;
            15'd4822: data <= 8'hFF;
            15'd4823: data <= 8'hFF;
            15'd4824: data <= 8'hFF;
            15'd4825: data <= 8'h80;
            15'd4826: data <= 8'h00;
            15'd4827: data <= 8'h00;
            15'd4828: data <= 8'h00;
            15'd4829: data <= 8'h00;
            15'd4830: data <= 8'h00;
            15'd4831: data <= 8'h00;
            15'd4832: data <= 8'h00;
            15'd4833: data <= 8'h00;
            15'd4834: data <= 8'h01;
            15'd4835: data <= 8'hFF;
            15'd4836: data <= 8'hFF;
            15'd4837: data <= 8'hFF;
            15'd4838: data <= 8'hFF;
            15'd4839: data <= 8'hFF;
            15'd4840: data <= 8'hFF;
            15'd4841: data <= 8'hFF;
            15'd4842: data <= 8'hE0;
            15'd4843: data <= 8'h00;
            15'd4844: data <= 8'h0F;
            15'd4845: data <= 8'hFF;
            15'd4846: data <= 8'hFE;
            15'd4847: data <= 8'h3F;
            15'd4848: data <= 8'hFF;
            15'd4849: data <= 8'hFF;
            15'd4850: data <= 8'hFF;
            15'd4851: data <= 8'hFF;
            15'd4852: data <= 8'hFF;
            15'd4853: data <= 8'hFF;
            15'd4854: data <= 8'hFF;
            15'd4855: data <= 8'h80;
            15'd4856: data <= 8'h00;
            15'd4857: data <= 8'h00;
            15'd4858: data <= 8'h00;
            15'd4859: data <= 8'h00;
            15'd4860: data <= 8'h00;
            15'd4861: data <= 8'h00;
            15'd4862: data <= 8'h00;
            15'd4863: data <= 8'h00;
            15'd4864: data <= 8'h01;
            15'd4865: data <= 8'hFF;
            15'd4866: data <= 8'hFF;
            15'd4867: data <= 8'hFF;
            15'd4868: data <= 8'hFF;
            15'd4869: data <= 8'hFF;
            15'd4870: data <= 8'hFF;
            15'd4871: data <= 8'hFF;
            15'd4872: data <= 8'hF7;
            15'd4873: data <= 8'hFF;
            15'd4874: data <= 8'hFF;
            15'd4875: data <= 8'hFF;
            15'd4876: data <= 8'hFF;
            15'd4877: data <= 8'hFF;
            15'd4878: data <= 8'hFF;
            15'd4879: data <= 8'hFF;
            15'd4880: data <= 8'hFF;
            15'd4881: data <= 8'hFF;
            15'd4882: data <= 8'hFF;
            15'd4883: data <= 8'hFF;
            15'd4884: data <= 8'hFF;
            15'd4885: data <= 8'h80;
            15'd4886: data <= 8'h00;
            15'd4887: data <= 8'h00;
            15'd4888: data <= 8'h00;
            15'd4889: data <= 8'h00;
            15'd4890: data <= 8'h00;
            15'd4891: data <= 8'h00;
            15'd4892: data <= 8'h00;
            15'd4893: data <= 8'h00;
            15'd4894: data <= 8'h01;
            15'd4895: data <= 8'hFF;
            15'd4896: data <= 8'hFF;
            15'd4897: data <= 8'hFF;
            15'd4898: data <= 8'hFF;
            15'd4899: data <= 8'hFF;
            15'd4900: data <= 8'hFF;
            15'd4901: data <= 8'hFF;
            15'd4902: data <= 8'hFF;
            15'd4903: data <= 8'hFF;
            15'd4904: data <= 8'hFF;
            15'd4905: data <= 8'hFF;
            15'd4906: data <= 8'hFF;
            15'd4907: data <= 8'hFF;
            15'd4908: data <= 8'hFF;
            15'd4909: data <= 8'hFF;
            15'd4910: data <= 8'hFF;
            15'd4911: data <= 8'hFF;
            15'd4912: data <= 8'hFF;
            15'd4913: data <= 8'hFF;
            15'd4914: data <= 8'hFF;
            15'd4915: data <= 8'h80;
            15'd4916: data <= 8'h00;
            15'd4917: data <= 8'h00;
            15'd4918: data <= 8'h00;
            15'd4919: data <= 8'h00;
            15'd4920: data <= 8'h00;
            15'd4921: data <= 8'h00;
            15'd4922: data <= 8'h00;
            15'd4923: data <= 8'h00;
            15'd4924: data <= 8'h01;
            15'd4925: data <= 8'hFF;
            15'd4926: data <= 8'hFF;
            15'd4927: data <= 8'hFF;
            15'd4928: data <= 8'hFF;
            15'd4929: data <= 8'hFF;
            15'd4930: data <= 8'hFF;
            15'd4931: data <= 8'hFF;
            15'd4932: data <= 8'hFF;
            15'd4933: data <= 8'hFF;
            15'd4934: data <= 8'hFF;
            15'd4935: data <= 8'hFF;
            15'd4936: data <= 8'hFF;
            15'd4937: data <= 8'hFF;
            15'd4938: data <= 8'hFF;
            15'd4939: data <= 8'hFF;
            15'd4940: data <= 8'hFF;
            15'd4941: data <= 8'hFF;
            15'd4942: data <= 8'hFF;
            15'd4943: data <= 8'hFF;
            15'd4944: data <= 8'hFF;
            15'd4945: data <= 8'h80;
            15'd4946: data <= 8'h00;
            15'd4947: data <= 8'h00;
            15'd4948: data <= 8'h00;
            15'd4949: data <= 8'h00;
            15'd4950: data <= 8'h00;
            15'd4951: data <= 8'h00;
            15'd4952: data <= 8'h00;
            15'd4953: data <= 8'h00;
            15'd4954: data <= 8'h01;
            15'd4955: data <= 8'hFF;
            15'd4956: data <= 8'hFF;
            15'd4957: data <= 8'hFF;
            15'd4958: data <= 8'hFF;
            15'd4959: data <= 8'hFF;
            15'd4960: data <= 8'hFF;
            15'd4961: data <= 8'hFF;
            15'd4962: data <= 8'hFF;
            15'd4963: data <= 8'hFF;
            15'd4964: data <= 8'hFF;
            15'd4965: data <= 8'hFF;
            15'd4966: data <= 8'hFF;
            15'd4967: data <= 8'hFF;
            15'd4968: data <= 8'hFF;
            15'd4969: data <= 8'hFF;
            15'd4970: data <= 8'hFF;
            15'd4971: data <= 8'hFF;
            15'd4972: data <= 8'hFF;
            15'd4973: data <= 8'hFF;
            15'd4974: data <= 8'hFF;
            15'd4975: data <= 8'h80;
            15'd4976: data <= 8'h00;
            15'd4977: data <= 8'h00;
            15'd4978: data <= 8'h00;
            15'd4979: data <= 8'h00;
            15'd4980: data <= 8'h00;
            15'd4981: data <= 8'h00;
            15'd4982: data <= 8'h00;
            15'd4983: data <= 8'h00;
            15'd4984: data <= 8'h01;
            15'd4985: data <= 8'hFF;
            15'd4986: data <= 8'hFF;
            15'd4987: data <= 8'hFF;
            15'd4988: data <= 8'hFF;
            15'd4989: data <= 8'hFF;
            15'd4990: data <= 8'hFF;
            15'd4991: data <= 8'hFF;
            15'd4992: data <= 8'hFF;
            15'd4993: data <= 8'hFF;
            15'd4994: data <= 8'hFF;
            15'd4995: data <= 8'hFF;
            15'd4996: data <= 8'hFF;
            15'd4997: data <= 8'hFF;
            15'd4998: data <= 8'hFF;
            15'd4999: data <= 8'hFF;
            15'd5000: data <= 8'hFF;
            15'd5001: data <= 8'hFF;
            15'd5002: data <= 8'hFF;
            15'd5003: data <= 8'hFF;
            15'd5004: data <= 8'hFF;
            15'd5005: data <= 8'h80;
            15'd5006: data <= 8'h00;
            15'd5007: data <= 8'h00;
            15'd5008: data <= 8'h00;
            15'd5009: data <= 8'h00;
            15'd5010: data <= 8'h00;
            15'd5011: data <= 8'h00;
            15'd5012: data <= 8'h00;
            15'd5013: data <= 8'h00;
            15'd5014: data <= 8'h01;
            15'd5015: data <= 8'hFF;
            15'd5016: data <= 8'hFF;
            15'd5017: data <= 8'hFF;
            15'd5018: data <= 8'hFF;
            15'd5019: data <= 8'hFF;
            15'd5020: data <= 8'hFF;
            15'd5021: data <= 8'hFF;
            15'd5022: data <= 8'hFF;
            15'd5023: data <= 8'hFF;
            15'd5024: data <= 8'hFF;
            15'd5025: data <= 8'hFF;
            15'd5026: data <= 8'hFF;
            15'd5027: data <= 8'hFF;
            15'd5028: data <= 8'hFF;
            15'd5029: data <= 8'hFF;
            15'd5030: data <= 8'hFF;
            15'd5031: data <= 8'hFF;
            15'd5032: data <= 8'hFF;
            15'd5033: data <= 8'hFF;
            15'd5034: data <= 8'hFF;
            15'd5035: data <= 8'h80;
            15'd5036: data <= 8'h00;
            15'd5037: data <= 8'h00;
            15'd5038: data <= 8'h00;
            15'd5039: data <= 8'h00;
            15'd5040: data <= 8'h00;
            15'd5041: data <= 8'h00;
            15'd5042: data <= 8'h00;
            15'd5043: data <= 8'h00;
            15'd5044: data <= 8'h01;
            15'd5045: data <= 8'hFF;
            15'd5046: data <= 8'hFF;
            15'd5047: data <= 8'hFF;
            15'd5048: data <= 8'hFF;
            15'd5049: data <= 8'hFF;
            15'd5050: data <= 8'hFF;
            15'd5051: data <= 8'hFF;
            15'd5052: data <= 8'hFF;
            15'd5053: data <= 8'hFF;
            15'd5054: data <= 8'hFF;
            15'd5055: data <= 8'hFF;
            15'd5056: data <= 8'hFF;
            15'd5057: data <= 8'hFF;
            15'd5058: data <= 8'hFF;
            15'd5059: data <= 8'hFF;
            15'd5060: data <= 8'hFF;
            15'd5061: data <= 8'hFF;
            15'd5062: data <= 8'hFF;
            15'd5063: data <= 8'hFF;
            15'd5064: data <= 8'hFF;
            15'd5065: data <= 8'h80;
            15'd5066: data <= 8'h00;
            15'd5067: data <= 8'h00;
            15'd5068: data <= 8'h00;
            15'd5069: data <= 8'h00;
            15'd5070: data <= 8'h00;
            15'd5071: data <= 8'h00;
            15'd5072: data <= 8'h00;
            15'd5073: data <= 8'h00;
            15'd5074: data <= 8'h01;
            15'd5075: data <= 8'hFF;
            15'd5076: data <= 8'hFF;
            15'd5077: data <= 8'hFF;
            15'd5078: data <= 8'hFF;
            15'd5079: data <= 8'hFF;
            15'd5080: data <= 8'hFF;
            15'd5081: data <= 8'hFF;
            15'd5082: data <= 8'hFF;
            15'd5083: data <= 8'hFF;
            15'd5084: data <= 8'hFF;
            15'd5085: data <= 8'hFF;
            15'd5086: data <= 8'hFF;
            15'd5087: data <= 8'hFF;
            15'd5088: data <= 8'hFF;
            15'd5089: data <= 8'hFF;
            15'd5090: data <= 8'hFF;
            15'd5091: data <= 8'hFF;
            15'd5092: data <= 8'hFF;
            15'd5093: data <= 8'hFF;
            15'd5094: data <= 8'hFF;
            15'd5095: data <= 8'h80;
            15'd5096: data <= 8'h00;
            15'd5097: data <= 8'h00;
            15'd5098: data <= 8'h00;
            15'd5099: data <= 8'h00;
            15'd5100: data <= 8'h00;
            15'd5101: data <= 8'h00;
            15'd5102: data <= 8'h00;
            15'd5103: data <= 8'h00;
            15'd5104: data <= 8'h01;
            15'd5105: data <= 8'hFF;
            15'd5106: data <= 8'hFF;
            15'd5107: data <= 8'hFF;
            15'd5108: data <= 8'hFF;
            15'd5109: data <= 8'hFF;
            15'd5110: data <= 8'hFF;
            15'd5111: data <= 8'hFF;
            15'd5112: data <= 8'hFF;
            15'd5113: data <= 8'hFF;
            15'd5114: data <= 8'hFF;
            15'd5115: data <= 8'hFF;
            15'd5116: data <= 8'hFF;
            15'd5117: data <= 8'hFF;
            15'd5118: data <= 8'hFF;
            15'd5119: data <= 8'hFF;
            15'd5120: data <= 8'hFF;
            15'd5121: data <= 8'hFF;
            15'd5122: data <= 8'hFF;
            15'd5123: data <= 8'hFF;
            15'd5124: data <= 8'hFF;
            15'd5125: data <= 8'h80;
            15'd5126: data <= 8'h00;
            15'd5127: data <= 8'h00;
            15'd5128: data <= 8'h00;
            15'd5129: data <= 8'h00;
            15'd5130: data <= 8'h00;
            15'd5131: data <= 8'h00;
            15'd5132: data <= 8'h00;
            15'd5133: data <= 8'h00;
            15'd5134: data <= 8'h01;
            15'd5135: data <= 8'hFF;
            15'd5136: data <= 8'hFF;
            15'd5137: data <= 8'hFF;
            15'd5138: data <= 8'hFF;
            15'd5139: data <= 8'hFF;
            15'd5140: data <= 8'hFF;
            15'd5141: data <= 8'hFF;
            15'd5142: data <= 8'hFF;
            15'd5143: data <= 8'hFF;
            15'd5144: data <= 8'hFF;
            15'd5145: data <= 8'hFF;
            15'd5146: data <= 8'hFF;
            15'd5147: data <= 8'hFF;
            15'd5148: data <= 8'hFF;
            15'd5149: data <= 8'hFF;
            15'd5150: data <= 8'hFF;
            15'd5151: data <= 8'hFF;
            15'd5152: data <= 8'hFF;
            15'd5153: data <= 8'hFF;
            15'd5154: data <= 8'hFF;
            15'd5155: data <= 8'h80;
            15'd5156: data <= 8'h00;
            15'd5157: data <= 8'h00;
            15'd5158: data <= 8'h00;
            15'd5159: data <= 8'h00;
            15'd5160: data <= 8'h00;
            15'd5161: data <= 8'h00;
            15'd5162: data <= 8'h00;
            15'd5163: data <= 8'h00;
            15'd5164: data <= 8'h01;
            15'd5165: data <= 8'hFF;
            15'd5166: data <= 8'hFF;
            15'd5167: data <= 8'hFF;
            15'd5168: data <= 8'hFF;
            15'd5169: data <= 8'hFF;
            15'd5170: data <= 8'hFF;
            15'd5171: data <= 8'hFF;
            15'd5172: data <= 8'hFF;
            15'd5173: data <= 8'hFF;
            15'd5174: data <= 8'hFF;
            15'd5175: data <= 8'hFF;
            15'd5176: data <= 8'hFF;
            15'd5177: data <= 8'hFF;
            15'd5178: data <= 8'hFF;
            15'd5179: data <= 8'hFF;
            15'd5180: data <= 8'hFF;
            15'd5181: data <= 8'hFF;
            15'd5182: data <= 8'hFF;
            15'd5183: data <= 8'hFF;
            15'd5184: data <= 8'hFF;
            15'd5185: data <= 8'h80;
            15'd5186: data <= 8'h00;
            15'd5187: data <= 8'h00;
            15'd5188: data <= 8'h00;
            15'd5189: data <= 8'h00;
            15'd5190: data <= 8'h00;
            15'd5191: data <= 8'h00;
            15'd5192: data <= 8'h00;
            15'd5193: data <= 8'h00;
            15'd5194: data <= 8'h01;
            15'd5195: data <= 8'hFF;
            15'd5196: data <= 8'hFF;
            15'd5197: data <= 8'hFF;
            15'd5198: data <= 8'hFF;
            15'd5199: data <= 8'hFF;
            15'd5200: data <= 8'hFF;
            15'd5201: data <= 8'hFF;
            15'd5202: data <= 8'hFF;
            15'd5203: data <= 8'hFF;
            15'd5204: data <= 8'hFF;
            15'd5205: data <= 8'hFF;
            15'd5206: data <= 8'hFF;
            15'd5207: data <= 8'hFF;
            15'd5208: data <= 8'hFF;
            15'd5209: data <= 8'hFF;
            15'd5210: data <= 8'hFF;
            15'd5211: data <= 8'hFF;
            15'd5212: data <= 8'hFF;
            15'd5213: data <= 8'hFF;
            15'd5214: data <= 8'hFF;
            15'd5215: data <= 8'h80;
            15'd5216: data <= 8'h00;
            15'd5217: data <= 8'h00;
            15'd5218: data <= 8'h00;
            15'd5219: data <= 8'h00;
            15'd5220: data <= 8'h00;
            15'd5221: data <= 8'h00;
            15'd5222: data <= 8'h00;
            15'd5223: data <= 8'h00;
            15'd5224: data <= 8'h01;
            15'd5225: data <= 8'hFF;
            15'd5226: data <= 8'hFF;
            15'd5227: data <= 8'hFF;
            15'd5228: data <= 8'hFF;
            15'd5229: data <= 8'hFF;
            15'd5230: data <= 8'hFF;
            15'd5231: data <= 8'hFF;
            15'd5232: data <= 8'hFF;
            15'd5233: data <= 8'hFF;
            15'd5234: data <= 8'hFF;
            15'd5235: data <= 8'hFF;
            15'd5236: data <= 8'hFF;
            15'd5237: data <= 8'hFF;
            15'd5238: data <= 8'hFF;
            15'd5239: data <= 8'hFF;
            15'd5240: data <= 8'hFF;
            15'd5241: data <= 8'hFF;
            15'd5242: data <= 8'hFF;
            15'd5243: data <= 8'hFF;
            15'd5244: data <= 8'hFF;
            15'd5245: data <= 8'h80;
            15'd5246: data <= 8'h00;
            15'd5247: data <= 8'h00;
            15'd5248: data <= 8'h00;
            15'd5249: data <= 8'h00;
            15'd5250: data <= 8'h00;
            15'd5251: data <= 8'h00;
            15'd5252: data <= 8'h00;
            15'd5253: data <= 8'h00;
            15'd5254: data <= 8'h01;
            15'd5255: data <= 8'hFF;
            15'd5256: data <= 8'hFF;
            15'd5257: data <= 8'hFF;
            15'd5258: data <= 8'hFF;
            15'd5259: data <= 8'hFF;
            15'd5260: data <= 8'hFF;
            15'd5261: data <= 8'hFF;
            15'd5262: data <= 8'hFF;
            15'd5263: data <= 8'hFF;
            15'd5264: data <= 8'hFF;
            15'd5265: data <= 8'hFF;
            15'd5266: data <= 8'hFF;
            15'd5267: data <= 8'hFF;
            15'd5268: data <= 8'hFF;
            15'd5269: data <= 8'hFF;
            15'd5270: data <= 8'hFF;
            15'd5271: data <= 8'hFF;
            15'd5272: data <= 8'hFF;
            15'd5273: data <= 8'hFF;
            15'd5274: data <= 8'hFF;
            15'd5275: data <= 8'h80;
            15'd5276: data <= 8'h00;
            15'd5277: data <= 8'h00;
            15'd5278: data <= 8'h00;
            15'd5279: data <= 8'h00;
            15'd5280: data <= 8'h00;
            15'd5281: data <= 8'h00;
            15'd5282: data <= 8'h00;
            15'd5283: data <= 8'h00;
            15'd5284: data <= 8'h01;
            15'd5285: data <= 8'hFF;
            15'd5286: data <= 8'hFF;
            15'd5287: data <= 8'hFF;
            15'd5288: data <= 8'hFF;
            15'd5289: data <= 8'hFF;
            15'd5290: data <= 8'hFF;
            15'd5291: data <= 8'hFF;
            15'd5292: data <= 8'hFF;
            15'd5293: data <= 8'hFF;
            15'd5294: data <= 8'hFF;
            15'd5295: data <= 8'hFF;
            15'd5296: data <= 8'hFF;
            15'd5297: data <= 8'hFF;
            15'd5298: data <= 8'hFF;
            15'd5299: data <= 8'hFF;
            15'd5300: data <= 8'hFF;
            15'd5301: data <= 8'hFF;
            15'd5302: data <= 8'hFF;
            15'd5303: data <= 8'hFF;
            15'd5304: data <= 8'hFF;
            15'd5305: data <= 8'h80;
            15'd5306: data <= 8'h00;
            15'd5307: data <= 8'h00;
            15'd5308: data <= 8'h00;
            15'd5309: data <= 8'h00;
            15'd5310: data <= 8'h00;
            15'd5311: data <= 8'h00;
            15'd5312: data <= 8'h00;
            15'd5313: data <= 8'h00;
            15'd5314: data <= 8'h01;
            15'd5315: data <= 8'hFF;
            15'd5316: data <= 8'hFF;
            15'd5317: data <= 8'hFF;
            15'd5318: data <= 8'hFF;
            15'd5319: data <= 8'hFF;
            15'd5320: data <= 8'hFF;
            15'd5321: data <= 8'hFF;
            15'd5322: data <= 8'hFF;
            15'd5323: data <= 8'hFF;
            15'd5324: data <= 8'hFF;
            15'd5325: data <= 8'hFF;
            15'd5326: data <= 8'hFF;
            15'd5327: data <= 8'hFF;
            15'd5328: data <= 8'hFF;
            15'd5329: data <= 8'hFF;
            15'd5330: data <= 8'hFF;
            15'd5331: data <= 8'hFF;
            15'd5332: data <= 8'hFF;
            15'd5333: data <= 8'hFF;
            15'd5334: data <= 8'hFF;
            15'd5335: data <= 8'h80;
            15'd5336: data <= 8'h00;
            15'd5337: data <= 8'h00;
            15'd5338: data <= 8'h00;
            15'd5339: data <= 8'h00;
            15'd5340: data <= 8'h00;
            15'd5341: data <= 8'h00;
            15'd5342: data <= 8'h00;
            15'd5343: data <= 8'h00;
            15'd5344: data <= 8'h01;
            15'd5345: data <= 8'hFF;
            15'd5346: data <= 8'hFF;
            15'd5347: data <= 8'hFF;
            15'd5348: data <= 8'hFF;
            15'd5349: data <= 8'hFF;
            15'd5350: data <= 8'hFF;
            15'd5351: data <= 8'hFF;
            15'd5352: data <= 8'hFF;
            15'd5353: data <= 8'hFF;
            15'd5354: data <= 8'hFF;
            15'd5355: data <= 8'hFF;
            15'd5356: data <= 8'hFF;
            15'd5357: data <= 8'hFF;
            15'd5358: data <= 8'hFF;
            15'd5359: data <= 8'hFF;
            15'd5360: data <= 8'hFF;
            15'd5361: data <= 8'hFF;
            15'd5362: data <= 8'hFF;
            15'd5363: data <= 8'hFF;
            15'd5364: data <= 8'hFF;
            15'd5365: data <= 8'h80;
            15'd5366: data <= 8'h00;
            15'd5367: data <= 8'h00;
            15'd5368: data <= 8'h00;
            15'd5369: data <= 8'h00;
            15'd5370: data <= 8'h00;
            15'd5371: data <= 8'h00;
            15'd5372: data <= 8'h00;
            15'd5373: data <= 8'h00;
            15'd5374: data <= 8'h01;
            15'd5375: data <= 8'hFF;
            15'd5376: data <= 8'hFF;
            15'd5377: data <= 8'hFF;
            15'd5378: data <= 8'hFF;
            15'd5379: data <= 8'hFF;
            15'd5380: data <= 8'hFF;
            15'd5381: data <= 8'hFF;
            15'd5382: data <= 8'hFF;
            15'd5383: data <= 8'hFF;
            15'd5384: data <= 8'hFF;
            15'd5385: data <= 8'hFF;
            15'd5386: data <= 8'hFF;
            15'd5387: data <= 8'hFF;
            15'd5388: data <= 8'hFF;
            15'd5389: data <= 8'hFF;
            15'd5390: data <= 8'hFF;
            15'd5391: data <= 8'hFF;
            15'd5392: data <= 8'hFF;
            15'd5393: data <= 8'hFF;
            15'd5394: data <= 8'hFF;
            15'd5395: data <= 8'h80;
            15'd5396: data <= 8'h00;
            15'd5397: data <= 8'h00;
            15'd5398: data <= 8'h00;
            15'd5399: data <= 8'h00;
            15'd5400: data <= 8'h00;
            15'd5401: data <= 8'h00;
            15'd5402: data <= 8'h00;
            15'd5403: data <= 8'h00;
            15'd5404: data <= 8'h01;
            15'd5405: data <= 8'hFF;
            15'd5406: data <= 8'hFF;
            15'd5407: data <= 8'hFF;
            15'd5408: data <= 8'hFF;
            15'd5409: data <= 8'hFF;
            15'd5410: data <= 8'hFF;
            15'd5411: data <= 8'hFF;
            15'd5412: data <= 8'hFF;
            15'd5413: data <= 8'hFF;
            15'd5414: data <= 8'hFF;
            15'd5415: data <= 8'hFF;
            15'd5416: data <= 8'hFF;
            15'd5417: data <= 8'hFF;
            15'd5418: data <= 8'hFF;
            15'd5419: data <= 8'hFF;
            15'd5420: data <= 8'hFF;
            15'd5421: data <= 8'hFF;
            15'd5422: data <= 8'hFF;
            15'd5423: data <= 8'hFF;
            15'd5424: data <= 8'hFF;
            15'd5425: data <= 8'h80;
            15'd5426: data <= 8'h00;
            15'd5427: data <= 8'h00;
            15'd5428: data <= 8'h00;
            15'd5429: data <= 8'h00;
            15'd5430: data <= 8'h00;
            15'd5431: data <= 8'h00;
            15'd5432: data <= 8'h00;
            15'd5433: data <= 8'h00;
            15'd5434: data <= 8'h01;
            15'd5435: data <= 8'hFF;
            15'd5436: data <= 8'hFF;
            15'd5437: data <= 8'hFF;
            15'd5438: data <= 8'hFF;
            15'd5439: data <= 8'hFF;
            15'd5440: data <= 8'hFF;
            15'd5441: data <= 8'hFF;
            15'd5442: data <= 8'hFF;
            15'd5443: data <= 8'hFF;
            15'd5444: data <= 8'hFF;
            15'd5445: data <= 8'hFF;
            15'd5446: data <= 8'hFF;
            15'd5447: data <= 8'hFF;
            15'd5448: data <= 8'hFF;
            15'd5449: data <= 8'hFF;
            15'd5450: data <= 8'hFF;
            15'd5451: data <= 8'hFF;
            15'd5452: data <= 8'hFF;
            15'd5453: data <= 8'hFF;
            15'd5454: data <= 8'hFF;
            15'd5455: data <= 8'h80;
            15'd5456: data <= 8'h00;
            15'd5457: data <= 8'h00;
            15'd5458: data <= 8'h00;
            15'd5459: data <= 8'h00;
            15'd5460: data <= 8'h00;
            15'd5461: data <= 8'h00;
            15'd5462: data <= 8'h00;
            15'd5463: data <= 8'h00;
            15'd5464: data <= 8'h01;
            15'd5465: data <= 8'hFF;
            15'd5466: data <= 8'hFF;
            15'd5467: data <= 8'hFF;
            15'd5468: data <= 8'hFF;
            15'd5469: data <= 8'hFF;
            15'd5470: data <= 8'hFF;
            15'd5471: data <= 8'hFF;
            15'd5472: data <= 8'hFF;
            15'd5473: data <= 8'hFF;
            15'd5474: data <= 8'hFF;
            15'd5475: data <= 8'hFF;
            15'd5476: data <= 8'hFF;
            15'd5477: data <= 8'hFF;
            15'd5478: data <= 8'hFF;
            15'd5479: data <= 8'hFF;
            15'd5480: data <= 8'hFF;
            15'd5481: data <= 8'hFF;
            15'd5482: data <= 8'hFF;
            15'd5483: data <= 8'hFF;
            15'd5484: data <= 8'hFF;
            15'd5485: data <= 8'h80;
            15'd5486: data <= 8'h00;
            15'd5487: data <= 8'h00;
            15'd5488: data <= 8'h00;
            15'd5489: data <= 8'h00;
            15'd5490: data <= 8'h00;
            15'd5491: data <= 8'h00;
            15'd5492: data <= 8'h00;
            15'd5493: data <= 8'h00;
            15'd5494: data <= 8'h01;
            15'd5495: data <= 8'hFF;
            15'd5496: data <= 8'hFF;
            15'd5497: data <= 8'hFF;
            15'd5498: data <= 8'hFF;
            15'd5499: data <= 8'hFF;
            15'd5500: data <= 8'hFF;
            15'd5501: data <= 8'hFF;
            15'd5502: data <= 8'hFF;
            15'd5503: data <= 8'hFF;
            15'd5504: data <= 8'hFF;
            15'd5505: data <= 8'hFF;
            15'd5506: data <= 8'hFF;
            15'd5507: data <= 8'hFF;
            15'd5508: data <= 8'hFF;
            15'd5509: data <= 8'hFF;
            15'd5510: data <= 8'hFF;
            15'd5511: data <= 8'hFF;
            15'd5512: data <= 8'hFF;
            15'd5513: data <= 8'hFF;
            15'd5514: data <= 8'hFF;
            15'd5515: data <= 8'h80;
            15'd5516: data <= 8'h00;
            15'd5517: data <= 8'h00;
            15'd5518: data <= 8'h00;
            15'd5519: data <= 8'h00;
            15'd5520: data <= 8'h00;
            15'd5521: data <= 8'h00;
            15'd5522: data <= 8'h00;
            15'd5523: data <= 8'h00;
            15'd5524: data <= 8'h01;
            15'd5525: data <= 8'hFF;
            15'd5526: data <= 8'hFF;
            15'd5527: data <= 8'hFF;
            15'd5528: data <= 8'hFF;
            15'd5529: data <= 8'hFF;
            15'd5530: data <= 8'hFF;
            15'd5531: data <= 8'hFF;
            15'd5532: data <= 8'hFF;
            15'd5533: data <= 8'hFF;
            15'd5534: data <= 8'hFF;
            15'd5535: data <= 8'hFF;
            15'd5536: data <= 8'hFF;
            15'd5537: data <= 8'hFF;
            15'd5538: data <= 8'hFF;
            15'd5539: data <= 8'hFF;
            15'd5540: data <= 8'hFF;
            15'd5541: data <= 8'hFF;
            15'd5542: data <= 8'hFF;
            15'd5543: data <= 8'hFF;
            15'd5544: data <= 8'hFF;
            15'd5545: data <= 8'h80;
            15'd5546: data <= 8'h00;
            15'd5547: data <= 8'h00;
            15'd5548: data <= 8'h00;
            15'd5549: data <= 8'h00;
            15'd5550: data <= 8'h00;
            15'd5551: data <= 8'h00;
            15'd5552: data <= 8'h00;
            15'd5553: data <= 8'h00;
            15'd5554: data <= 8'h01;
            15'd5555: data <= 8'hFF;
            15'd5556: data <= 8'hFF;
            15'd5557: data <= 8'hFF;
            15'd5558: data <= 8'hFF;
            15'd5559: data <= 8'hFF;
            15'd5560: data <= 8'hFF;
            15'd5561: data <= 8'hFF;
            15'd5562: data <= 8'hFF;
            15'd5563: data <= 8'hFF;
            15'd5564: data <= 8'hFF;
            15'd5565: data <= 8'hFF;
            15'd5566: data <= 8'hFF;
            15'd5567: data <= 8'hFF;
            15'd5568: data <= 8'hFF;
            15'd5569: data <= 8'hFF;
            15'd5570: data <= 8'hFF;
            15'd5571: data <= 8'hFF;
            15'd5572: data <= 8'hFF;
            15'd5573: data <= 8'hFF;
            15'd5574: data <= 8'hFF;
            15'd5575: data <= 8'h80;
            15'd5576: data <= 8'h00;
            15'd5577: data <= 8'h00;
            15'd5578: data <= 8'h00;
            15'd5579: data <= 8'h00;
            15'd5580: data <= 8'h00;
            15'd5581: data <= 8'h00;
            15'd5582: data <= 8'h00;
            15'd5583: data <= 8'h00;
            15'd5584: data <= 8'h01;
            15'd5585: data <= 8'hFF;
            15'd5586: data <= 8'hFF;
            15'd5587: data <= 8'hFF;
            15'd5588: data <= 8'hFF;
            15'd5589: data <= 8'hFF;
            15'd5590: data <= 8'hFF;
            15'd5591: data <= 8'hFF;
            15'd5592: data <= 8'hFF;
            15'd5593: data <= 8'hFF;
            15'd5594: data <= 8'hFF;
            15'd5595: data <= 8'hFF;
            15'd5596: data <= 8'hFF;
            15'd5597: data <= 8'hFF;
            15'd5598: data <= 8'hFF;
            15'd5599: data <= 8'hFF;
            15'd5600: data <= 8'hFF;
            15'd5601: data <= 8'hFF;
            15'd5602: data <= 8'hFF;
            15'd5603: data <= 8'hFF;
            15'd5604: data <= 8'hFF;
            15'd5605: data <= 8'h80;
            15'd5606: data <= 8'h00;
            15'd5607: data <= 8'h00;
            15'd5608: data <= 8'h00;
            15'd5609: data <= 8'h00;
            15'd5610: data <= 8'h00;
            15'd5611: data <= 8'h00;
            15'd5612: data <= 8'h00;
            15'd5613: data <= 8'h00;
            15'd5614: data <= 8'h01;
            15'd5615: data <= 8'hFF;
            15'd5616: data <= 8'hFF;
            15'd5617: data <= 8'hFF;
            15'd5618: data <= 8'hFF;
            15'd5619: data <= 8'hFF;
            15'd5620: data <= 8'hFF;
            15'd5621: data <= 8'hFF;
            15'd5622: data <= 8'hFF;
            15'd5623: data <= 8'hFF;
            15'd5624: data <= 8'hFF;
            15'd5625: data <= 8'hFF;
            15'd5626: data <= 8'hFF;
            15'd5627: data <= 8'hFF;
            15'd5628: data <= 8'hFF;
            15'd5629: data <= 8'hFF;
            15'd5630: data <= 8'hFF;
            15'd5631: data <= 8'hFF;
            15'd5632: data <= 8'hFF;
            15'd5633: data <= 8'hFF;
            15'd5634: data <= 8'hFF;
            15'd5635: data <= 8'h80;
            15'd5636: data <= 8'h00;
            15'd5637: data <= 8'h00;
            15'd5638: data <= 8'h00;
            15'd5639: data <= 8'h00;
            15'd5640: data <= 8'h00;
            15'd5641: data <= 8'h00;
            15'd5642: data <= 8'h00;
            15'd5643: data <= 8'h00;
            15'd5644: data <= 8'h01;
            15'd5645: data <= 8'hFF;
            15'd5646: data <= 8'hFF;
            15'd5647: data <= 8'hFF;
            15'd5648: data <= 8'hFF;
            15'd5649: data <= 8'hFF;
            15'd5650: data <= 8'hFF;
            15'd5651: data <= 8'hFF;
            15'd5652: data <= 8'hFF;
            15'd5653: data <= 8'hFF;
            15'd5654: data <= 8'hFF;
            15'd5655: data <= 8'hFF;
            15'd5656: data <= 8'hFF;
            15'd5657: data <= 8'hFF;
            15'd5658: data <= 8'hFF;
            15'd5659: data <= 8'hFF;
            15'd5660: data <= 8'hFF;
            15'd5661: data <= 8'hFF;
            15'd5662: data <= 8'hFF;
            15'd5663: data <= 8'hFF;
            15'd5664: data <= 8'hFF;
            15'd5665: data <= 8'h80;
            15'd5666: data <= 8'h00;
            15'd5667: data <= 8'h00;
            15'd5668: data <= 8'h00;
            15'd5669: data <= 8'h00;
            15'd5670: data <= 8'h00;
            15'd5671: data <= 8'h00;
            15'd5672: data <= 8'h00;
            15'd5673: data <= 8'h00;
            15'd5674: data <= 8'h01;
            15'd5675: data <= 8'hFF;
            15'd5676: data <= 8'hFF;
            15'd5677: data <= 8'hFF;
            15'd5678: data <= 8'hFF;
            15'd5679: data <= 8'hFF;
            15'd5680: data <= 8'hFF;
            15'd5681: data <= 8'hFF;
            15'd5682: data <= 8'hFF;
            15'd5683: data <= 8'hFF;
            15'd5684: data <= 8'hFF;
            15'd5685: data <= 8'hFF;
            15'd5686: data <= 8'hFF;
            15'd5687: data <= 8'hFF;
            15'd5688: data <= 8'hFF;
            15'd5689: data <= 8'hFF;
            15'd5690: data <= 8'hFF;
            15'd5691: data <= 8'hFF;
            15'd5692: data <= 8'hFF;
            15'd5693: data <= 8'hFF;
            15'd5694: data <= 8'hFF;
            15'd5695: data <= 8'h80;
            15'd5696: data <= 8'h00;
            15'd5697: data <= 8'h00;
            15'd5698: data <= 8'h00;
            15'd5699: data <= 8'h00;
            15'd5700: data <= 8'h00;
            15'd5701: data <= 8'h00;
            15'd5702: data <= 8'h00;
            15'd5703: data <= 8'h00;
            15'd5704: data <= 8'h01;
            15'd5705: data <= 8'hFF;
            15'd5706: data <= 8'hFF;
            15'd5707: data <= 8'hFF;
            15'd5708: data <= 8'hFF;
            15'd5709: data <= 8'hFF;
            15'd5710: data <= 8'hFF;
            15'd5711: data <= 8'hFF;
            15'd5712: data <= 8'hFF;
            15'd5713: data <= 8'hFF;
            15'd5714: data <= 8'hFF;
            15'd5715: data <= 8'hFF;
            15'd5716: data <= 8'hFF;
            15'd5717: data <= 8'hFF;
            15'd5718: data <= 8'hFF;
            15'd5719: data <= 8'hFF;
            15'd5720: data <= 8'hFF;
            15'd5721: data <= 8'hFF;
            15'd5722: data <= 8'hFF;
            15'd5723: data <= 8'hFF;
            15'd5724: data <= 8'hFF;
            15'd5725: data <= 8'h80;
            15'd5726: data <= 8'h00;
            15'd5727: data <= 8'h00;
            15'd5728: data <= 8'h00;
            15'd5729: data <= 8'h00;
            15'd5730: data <= 8'h00;
            15'd5731: data <= 8'h00;
            15'd5732: data <= 8'h00;
            15'd5733: data <= 8'h00;
            15'd5734: data <= 8'h01;
            15'd5735: data <= 8'hFF;
            15'd5736: data <= 8'hFF;
            15'd5737: data <= 8'hFF;
            15'd5738: data <= 8'hFF;
            15'd5739: data <= 8'hFF;
            15'd5740: data <= 8'hFF;
            15'd5741: data <= 8'hFF;
            15'd5742: data <= 8'hFF;
            15'd5743: data <= 8'hFF;
            15'd5744: data <= 8'hFF;
            15'd5745: data <= 8'hFF;
            15'd5746: data <= 8'hFF;
            15'd5747: data <= 8'hFF;
            15'd5748: data <= 8'hFF;
            15'd5749: data <= 8'hFF;
            15'd5750: data <= 8'hFF;
            15'd5751: data <= 8'hFF;
            15'd5752: data <= 8'hFF;
            15'd5753: data <= 8'hFF;
            15'd5754: data <= 8'hFF;
            15'd5755: data <= 8'h80;
            15'd5756: data <= 8'h00;
            15'd5757: data <= 8'h00;
            15'd5758: data <= 8'h00;
            15'd5759: data <= 8'h00;
            15'd5760: data <= 8'h00;
            15'd5761: data <= 8'h00;
            15'd5762: data <= 8'h00;
            15'd5763: data <= 8'h00;
            15'd5764: data <= 8'h01;
            15'd5765: data <= 8'hFF;
            15'd5766: data <= 8'hFF;
            15'd5767: data <= 8'hFF;
            15'd5768: data <= 8'hFF;
            15'd5769: data <= 8'hFF;
            15'd5770: data <= 8'hFF;
            15'd5771: data <= 8'hFF;
            15'd5772: data <= 8'hFF;
            15'd5773: data <= 8'hFF;
            15'd5774: data <= 8'hFF;
            15'd5775: data <= 8'hFF;
            15'd5776: data <= 8'hFF;
            15'd5777: data <= 8'hFF;
            15'd5778: data <= 8'hFF;
            15'd5779: data <= 8'hFF;
            15'd5780: data <= 8'hFF;
            15'd5781: data <= 8'hFF;
            15'd5782: data <= 8'hFF;
            15'd5783: data <= 8'hFF;
            15'd5784: data <= 8'hFF;
            15'd5785: data <= 8'h80;
            15'd5786: data <= 8'h00;
            15'd5787: data <= 8'h00;
            15'd5788: data <= 8'h00;
            15'd5789: data <= 8'h00;
            15'd5790: data <= 8'h00;
            15'd5791: data <= 8'h00;
            15'd5792: data <= 8'h00;
            15'd5793: data <= 8'h00;
            15'd5794: data <= 8'h01;
            15'd5795: data <= 8'hFF;
            15'd5796: data <= 8'hFF;
            15'd5797: data <= 8'hFF;
            15'd5798: data <= 8'hFF;
            15'd5799: data <= 8'hFF;
            15'd5800: data <= 8'hFF;
            15'd5801: data <= 8'hFF;
            15'd5802: data <= 8'hFF;
            15'd5803: data <= 8'hFF;
            15'd5804: data <= 8'hFF;
            15'd5805: data <= 8'hFF;
            15'd5806: data <= 8'hFF;
            15'd5807: data <= 8'hFF;
            15'd5808: data <= 8'hFF;
            15'd5809: data <= 8'hFF;
            15'd5810: data <= 8'hFF;
            15'd5811: data <= 8'hFF;
            15'd5812: data <= 8'hFF;
            15'd5813: data <= 8'hFF;
            15'd5814: data <= 8'hFF;
            15'd5815: data <= 8'h80;
            15'd5816: data <= 8'h00;
            15'd5817: data <= 8'h00;
            15'd5818: data <= 8'h00;
            15'd5819: data <= 8'h00;
            15'd5820: data <= 8'h00;
            15'd5821: data <= 8'h00;
            15'd5822: data <= 8'h00;
            15'd5823: data <= 8'h00;
            15'd5824: data <= 8'h01;
            15'd5825: data <= 8'hFF;
            15'd5826: data <= 8'hFF;
            15'd5827: data <= 8'hFF;
            15'd5828: data <= 8'hFF;
            15'd5829: data <= 8'hFF;
            15'd5830: data <= 8'hFF;
            15'd5831: data <= 8'hFF;
            15'd5832: data <= 8'hFF;
            15'd5833: data <= 8'hFF;
            15'd5834: data <= 8'hFF;
            15'd5835: data <= 8'hFF;
            15'd5836: data <= 8'hFF;
            15'd5837: data <= 8'hFF;
            15'd5838: data <= 8'hFF;
            15'd5839: data <= 8'hFF;
            15'd5840: data <= 8'hFF;
            15'd5841: data <= 8'hFF;
            15'd5842: data <= 8'hFF;
            15'd5843: data <= 8'hFF;
            15'd5844: data <= 8'hFF;
            15'd5845: data <= 8'h80;
            15'd5846: data <= 8'h00;
            15'd5847: data <= 8'h00;
            15'd5848: data <= 8'h00;
            15'd5849: data <= 8'h00;
            15'd5850: data <= 8'h00;
            15'd5851: data <= 8'h00;
            15'd5852: data <= 8'h00;
            15'd5853: data <= 8'h00;
            15'd5854: data <= 8'h01;
            15'd5855: data <= 8'hFF;
            15'd5856: data <= 8'hFF;
            15'd5857: data <= 8'hFF;
            15'd5858: data <= 8'hFF;
            15'd5859: data <= 8'hFF;
            15'd5860: data <= 8'hFF;
            15'd5861: data <= 8'hFF;
            15'd5862: data <= 8'hFF;
            15'd5863: data <= 8'hFF;
            15'd5864: data <= 8'hFF;
            15'd5865: data <= 8'hFF;
            15'd5866: data <= 8'hFF;
            15'd5867: data <= 8'hFF;
            15'd5868: data <= 8'hFF;
            15'd5869: data <= 8'hFF;
            15'd5870: data <= 8'hFF;
            15'd5871: data <= 8'hFF;
            15'd5872: data <= 8'hFF;
            15'd5873: data <= 8'hFF;
            15'd5874: data <= 8'hFF;
            15'd5875: data <= 8'h80;
            15'd5876: data <= 8'h00;
            15'd5877: data <= 8'h00;
            15'd5878: data <= 8'h00;
            15'd5879: data <= 8'h00;
            15'd5880: data <= 8'h00;
            15'd5881: data <= 8'h00;
            15'd5882: data <= 8'h00;
            15'd5883: data <= 8'h00;
            15'd5884: data <= 8'h01;
            15'd5885: data <= 8'hFF;
            15'd5886: data <= 8'hFF;
            15'd5887: data <= 8'hFF;
            15'd5888: data <= 8'hFF;
            15'd5889: data <= 8'hFF;
            15'd5890: data <= 8'hFF;
            15'd5891: data <= 8'hFF;
            15'd5892: data <= 8'hFF;
            15'd5893: data <= 8'hFF;
            15'd5894: data <= 8'hFF;
            15'd5895: data <= 8'hFF;
            15'd5896: data <= 8'hFF;
            15'd5897: data <= 8'hFF;
            15'd5898: data <= 8'hFF;
            15'd5899: data <= 8'hFF;
            15'd5900: data <= 8'hFF;
            15'd5901: data <= 8'hFF;
            15'd5902: data <= 8'hFF;
            15'd5903: data <= 8'hFF;
            15'd5904: data <= 8'hFF;
            15'd5905: data <= 8'h80;
            15'd5906: data <= 8'h00;
            15'd5907: data <= 8'h00;
            15'd5908: data <= 8'h00;
            15'd5909: data <= 8'h00;
            15'd5910: data <= 8'h00;
            15'd5911: data <= 8'h00;
            15'd5912: data <= 8'h00;
            15'd5913: data <= 8'h00;
            15'd5914: data <= 8'h01;
            15'd5915: data <= 8'hFF;
            15'd5916: data <= 8'hFF;
            15'd5917: data <= 8'hFF;
            15'd5918: data <= 8'hFF;
            15'd5919: data <= 8'hFF;
            15'd5920: data <= 8'hFF;
            15'd5921: data <= 8'hFF;
            15'd5922: data <= 8'hFF;
            15'd5923: data <= 8'hFF;
            15'd5924: data <= 8'hFF;
            15'd5925: data <= 8'hFF;
            15'd5926: data <= 8'hFF;
            15'd5927: data <= 8'hFF;
            15'd5928: data <= 8'hFF;
            15'd5929: data <= 8'hFF;
            15'd5930: data <= 8'hFF;
            15'd5931: data <= 8'hFF;
            15'd5932: data <= 8'hFF;
            15'd5933: data <= 8'hFF;
            15'd5934: data <= 8'hFF;
            15'd5935: data <= 8'h80;
            15'd5936: data <= 8'h00;
            15'd5937: data <= 8'h00;
            15'd5938: data <= 8'h00;
            15'd5939: data <= 8'h00;
            15'd5940: data <= 8'h00;
            15'd5941: data <= 8'h00;
            15'd5942: data <= 8'h00;
            15'd5943: data <= 8'h00;
            15'd5944: data <= 8'h01;
            15'd5945: data <= 8'hFF;
            15'd5946: data <= 8'hFF;
            15'd5947: data <= 8'hFF;
            15'd5948: data <= 8'hFF;
            15'd5949: data <= 8'hFF;
            15'd5950: data <= 8'hFF;
            15'd5951: data <= 8'hFF;
            15'd5952: data <= 8'hFF;
            15'd5953: data <= 8'hFF;
            15'd5954: data <= 8'hFF;
            15'd5955: data <= 8'hFF;
            15'd5956: data <= 8'hFF;
            15'd5957: data <= 8'hFF;
            15'd5958: data <= 8'hFF;
            15'd5959: data <= 8'hFF;
            15'd5960: data <= 8'hFF;
            15'd5961: data <= 8'hFF;
            15'd5962: data <= 8'hFF;
            15'd5963: data <= 8'hFF;
            15'd5964: data <= 8'hFF;
            15'd5965: data <= 8'h80;
            15'd5966: data <= 8'h00;
            15'd5967: data <= 8'h00;
            15'd5968: data <= 8'h00;
            15'd5969: data <= 8'h00;
            15'd5970: data <= 8'h00;
            15'd5971: data <= 8'h00;
            15'd5972: data <= 8'h00;
            15'd5973: data <= 8'h00;
            15'd5974: data <= 8'h01;
            15'd5975: data <= 8'hFF;
            15'd5976: data <= 8'hFF;
            15'd5977: data <= 8'hFF;
            15'd5978: data <= 8'hFF;
            15'd5979: data <= 8'hFF;
            15'd5980: data <= 8'hFF;
            15'd5981: data <= 8'hFF;
            15'd5982: data <= 8'hFF;
            15'd5983: data <= 8'hFF;
            15'd5984: data <= 8'hFF;
            15'd5985: data <= 8'hFF;
            15'd5986: data <= 8'hFF;
            15'd5987: data <= 8'hFF;
            15'd5988: data <= 8'hFF;
            15'd5989: data <= 8'hFF;
            15'd5990: data <= 8'hFF;
            15'd5991: data <= 8'hFF;
            15'd5992: data <= 8'hFF;
            15'd5993: data <= 8'hFF;
            15'd5994: data <= 8'hFF;
            15'd5995: data <= 8'h80;
            15'd5996: data <= 8'h00;
            15'd5997: data <= 8'h00;
            15'd5998: data <= 8'h00;
            15'd5999: data <= 8'h00;
            15'd6000: data <= 8'h00;
            15'd6001: data <= 8'h00;
            15'd6002: data <= 8'h00;
            15'd6003: data <= 8'h00;
            15'd6004: data <= 8'h01;
            15'd6005: data <= 8'hFF;
            15'd6006: data <= 8'hFF;
            15'd6007: data <= 8'hFF;
            15'd6008: data <= 8'hFF;
            15'd6009: data <= 8'hFF;
            15'd6010: data <= 8'hFF;
            15'd6011: data <= 8'hFF;
            15'd6012: data <= 8'hFF;
            15'd6013: data <= 8'hFF;
            15'd6014: data <= 8'hFF;
            15'd6015: data <= 8'hFF;
            15'd6016: data <= 8'hFF;
            15'd6017: data <= 8'hFF;
            15'd6018: data <= 8'hFF;
            15'd6019: data <= 8'hFF;
            15'd6020: data <= 8'hFF;
            15'd6021: data <= 8'hFF;
            15'd6022: data <= 8'hFF;
            15'd6023: data <= 8'hFF;
            15'd6024: data <= 8'hFF;
            15'd6025: data <= 8'h80;
            15'd6026: data <= 8'h00;
            15'd6027: data <= 8'h00;
            15'd6028: data <= 8'h00;
            15'd6029: data <= 8'h00;
            15'd6030: data <= 8'h00;
            15'd6031: data <= 8'h00;
            15'd6032: data <= 8'h00;
            15'd6033: data <= 8'h00;
            15'd6034: data <= 8'h01;
            15'd6035: data <= 8'hFF;
            15'd6036: data <= 8'hFF;
            15'd6037: data <= 8'hFF;
            15'd6038: data <= 8'hFF;
            15'd6039: data <= 8'hFF;
            15'd6040: data <= 8'hFF;
            15'd6041: data <= 8'hFF;
            15'd6042: data <= 8'hFF;
            15'd6043: data <= 8'hFF;
            15'd6044: data <= 8'hFF;
            15'd6045: data <= 8'hFF;
            15'd6046: data <= 8'hFF;
            15'd6047: data <= 8'hFF;
            15'd6048: data <= 8'hFF;
            15'd6049: data <= 8'hFF;
            15'd6050: data <= 8'hFF;
            15'd6051: data <= 8'hFF;
            15'd6052: data <= 8'hFF;
            15'd6053: data <= 8'hFF;
            15'd6054: data <= 8'hFF;
            15'd6055: data <= 8'h80;
            15'd6056: data <= 8'h00;
            15'd6057: data <= 8'h00;
            15'd6058: data <= 8'h00;
            15'd6059: data <= 8'h00;
            15'd6060: data <= 8'h00;
            15'd6061: data <= 8'h00;
            15'd6062: data <= 8'h00;
            15'd6063: data <= 8'h00;
            15'd6064: data <= 8'h01;
            15'd6065: data <= 8'hFF;
            15'd6066: data <= 8'hFF;
            15'd6067: data <= 8'hFF;
            15'd6068: data <= 8'hFF;
            15'd6069: data <= 8'hFF;
            15'd6070: data <= 8'hFF;
            15'd6071: data <= 8'hFF;
            15'd6072: data <= 8'hFF;
            15'd6073: data <= 8'hFF;
            15'd6074: data <= 8'hFF;
            15'd6075: data <= 8'hFF;
            15'd6076: data <= 8'hFF;
            15'd6077: data <= 8'hFF;
            15'd6078: data <= 8'hFF;
            15'd6079: data <= 8'hFF;
            15'd6080: data <= 8'hFF;
            15'd6081: data <= 8'hFF;
            15'd6082: data <= 8'hFF;
            15'd6083: data <= 8'hFF;
            15'd6084: data <= 8'hFF;
            15'd6085: data <= 8'h80;
            15'd6086: data <= 8'h00;
            15'd6087: data <= 8'h00;
            15'd6088: data <= 8'h00;
            15'd6089: data <= 8'h00;
            15'd6090: data <= 8'h00;
            15'd6091: data <= 8'h00;
            15'd6092: data <= 8'h00;
            15'd6093: data <= 8'h00;
            15'd6094: data <= 8'h01;
            15'd6095: data <= 8'hFF;
            15'd6096: data <= 8'hFF;
            15'd6097: data <= 8'hFF;
            15'd6098: data <= 8'hFF;
            15'd6099: data <= 8'hFF;
            15'd6100: data <= 8'hFF;
            15'd6101: data <= 8'hFF;
            15'd6102: data <= 8'hFF;
            15'd6103: data <= 8'hFF;
            15'd6104: data <= 8'hFF;
            15'd6105: data <= 8'hFF;
            15'd6106: data <= 8'hFF;
            15'd6107: data <= 8'hFF;
            15'd6108: data <= 8'hFF;
            15'd6109: data <= 8'hFF;
            15'd6110: data <= 8'hFF;
            15'd6111: data <= 8'hFF;
            15'd6112: data <= 8'hFF;
            15'd6113: data <= 8'hFF;
            15'd6114: data <= 8'hFF;
            15'd6115: data <= 8'h80;
            15'd6116: data <= 8'h00;
            15'd6117: data <= 8'h00;
            15'd6118: data <= 8'h00;
            15'd6119: data <= 8'h00;
            15'd6120: data <= 8'h00;
            15'd6121: data <= 8'h00;
            15'd6122: data <= 8'h00;
            15'd6123: data <= 8'h00;
            15'd6124: data <= 8'h01;
            15'd6125: data <= 8'hFF;
            15'd6126: data <= 8'hFF;
            15'd6127: data <= 8'hFF;
            15'd6128: data <= 8'hFF;
            15'd6129: data <= 8'hFF;
            15'd6130: data <= 8'hFF;
            15'd6131: data <= 8'hFF;
            15'd6132: data <= 8'hFF;
            15'd6133: data <= 8'hFF;
            15'd6134: data <= 8'hFF;
            15'd6135: data <= 8'hFF;
            15'd6136: data <= 8'hFF;
            15'd6137: data <= 8'hFF;
            15'd6138: data <= 8'hFF;
            15'd6139: data <= 8'hFF;
            15'd6140: data <= 8'hFF;
            15'd6141: data <= 8'hFF;
            15'd6142: data <= 8'hFF;
            15'd6143: data <= 8'hFF;
            15'd6144: data <= 8'hFF;
            15'd6145: data <= 8'h80;
            15'd6146: data <= 8'h00;
            15'd6147: data <= 8'h00;
            15'd6148: data <= 8'h00;
            15'd6149: data <= 8'h00;
            15'd6150: data <= 8'h00;
            15'd6151: data <= 8'h00;
            15'd6152: data <= 8'h00;
            15'd6153: data <= 8'h00;
            15'd6154: data <= 8'h01;
            15'd6155: data <= 8'hFF;
            15'd6156: data <= 8'hFF;
            15'd6157: data <= 8'hFF;
            15'd6158: data <= 8'hFF;
            15'd6159: data <= 8'hFF;
            15'd6160: data <= 8'hFF;
            15'd6161: data <= 8'hFF;
            15'd6162: data <= 8'hFF;
            15'd6163: data <= 8'hFF;
            15'd6164: data <= 8'hFF;
            15'd6165: data <= 8'hFF;
            15'd6166: data <= 8'hFF;
            15'd6167: data <= 8'hFF;
            15'd6168: data <= 8'hFF;
            15'd6169: data <= 8'hFF;
            15'd6170: data <= 8'hFF;
            15'd6171: data <= 8'hFF;
            15'd6172: data <= 8'hFF;
            15'd6173: data <= 8'hFF;
            15'd6174: data <= 8'hFF;
            15'd6175: data <= 8'h80;
            15'd6176: data <= 8'h00;
            15'd6177: data <= 8'h00;
            15'd6178: data <= 8'h00;
            15'd6179: data <= 8'h00;
            15'd6180: data <= 8'h00;
            15'd6181: data <= 8'h00;
            15'd6182: data <= 8'h00;
            15'd6183: data <= 8'h00;
            15'd6184: data <= 8'h01;
            15'd6185: data <= 8'hFF;
            15'd6186: data <= 8'hFF;
            15'd6187: data <= 8'hFF;
            15'd6188: data <= 8'hFF;
            15'd6189: data <= 8'hFF;
            15'd6190: data <= 8'hFF;
            15'd6191: data <= 8'hFF;
            15'd6192: data <= 8'hFF;
            15'd6193: data <= 8'hFF;
            15'd6194: data <= 8'hFF;
            15'd6195: data <= 8'hFF;
            15'd6196: data <= 8'hFF;
            15'd6197: data <= 8'hFF;
            15'd6198: data <= 8'hFF;
            15'd6199: data <= 8'hFF;
            15'd6200: data <= 8'hFF;
            15'd6201: data <= 8'hFF;
            15'd6202: data <= 8'hFF;
            15'd6203: data <= 8'hFF;
            15'd6204: data <= 8'hFF;
            15'd6205: data <= 8'h80;
            15'd6206: data <= 8'h00;
            15'd6207: data <= 8'h00;
            15'd6208: data <= 8'h00;
            15'd6209: data <= 8'h00;
            15'd6210: data <= 8'h00;
            15'd6211: data <= 8'h00;
            15'd6212: data <= 8'h00;
            15'd6213: data <= 8'h00;
            15'd6214: data <= 8'h01;
            15'd6215: data <= 8'hFF;
            15'd6216: data <= 8'hFF;
            15'd6217: data <= 8'hFF;
            15'd6218: data <= 8'hFF;
            15'd6219: data <= 8'hFF;
            15'd6220: data <= 8'hFF;
            15'd6221: data <= 8'hFF;
            15'd6222: data <= 8'hFF;
            15'd6223: data <= 8'hFF;
            15'd6224: data <= 8'hFF;
            15'd6225: data <= 8'hFF;
            15'd6226: data <= 8'hFF;
            15'd6227: data <= 8'hFF;
            15'd6228: data <= 8'hFF;
            15'd6229: data <= 8'hFF;
            15'd6230: data <= 8'hFF;
            15'd6231: data <= 8'hFF;
            15'd6232: data <= 8'hFF;
            15'd6233: data <= 8'hFF;
            15'd6234: data <= 8'hFF;
            15'd6235: data <= 8'h80;
            15'd6236: data <= 8'h00;
            15'd6237: data <= 8'h00;
            15'd6238: data <= 8'h00;
            15'd6239: data <= 8'h00;
            15'd6240: data <= 8'h00;
            15'd6241: data <= 8'h00;
            15'd6242: data <= 8'h00;
            15'd6243: data <= 8'h00;
            15'd6244: data <= 8'h01;
            15'd6245: data <= 8'hFF;
            15'd6246: data <= 8'hFF;
            15'd6247: data <= 8'hFF;
            15'd6248: data <= 8'hFF;
            15'd6249: data <= 8'hFF;
            15'd6250: data <= 8'hFF;
            15'd6251: data <= 8'hFF;
            15'd6252: data <= 8'hFF;
            15'd6253: data <= 8'hFF;
            15'd6254: data <= 8'hFF;
            15'd6255: data <= 8'hFF;
            15'd6256: data <= 8'hFF;
            15'd6257: data <= 8'hFF;
            15'd6258: data <= 8'hFF;
            15'd6259: data <= 8'hFF;
            15'd6260: data <= 8'hFF;
            15'd6261: data <= 8'hFF;
            15'd6262: data <= 8'hFF;
            15'd6263: data <= 8'hFF;
            15'd6264: data <= 8'hFF;
            15'd6265: data <= 8'h80;
            15'd6266: data <= 8'h00;
            15'd6267: data <= 8'h00;
            15'd6268: data <= 8'h00;
            15'd6269: data <= 8'h00;
            15'd6270: data <= 8'h00;
            15'd6271: data <= 8'h00;
            15'd6272: data <= 8'h00;
            15'd6273: data <= 8'h00;
            15'd6274: data <= 8'h01;
            15'd6275: data <= 8'hFF;
            15'd6276: data <= 8'hFF;
            15'd6277: data <= 8'hFF;
            15'd6278: data <= 8'hFF;
            15'd6279: data <= 8'hFF;
            15'd6280: data <= 8'hFF;
            15'd6281: data <= 8'hFF;
            15'd6282: data <= 8'hFF;
            15'd6283: data <= 8'hFF;
            15'd6284: data <= 8'hFF;
            15'd6285: data <= 8'hFF;
            15'd6286: data <= 8'hFF;
            15'd6287: data <= 8'hFF;
            15'd6288: data <= 8'hFF;
            15'd6289: data <= 8'hFF;
            15'd6290: data <= 8'hFF;
            15'd6291: data <= 8'hFF;
            15'd6292: data <= 8'hFF;
            15'd6293: data <= 8'hFF;
            15'd6294: data <= 8'hFF;
            15'd6295: data <= 8'h80;
            15'd6296: data <= 8'h00;
            15'd6297: data <= 8'h00;
            15'd6298: data <= 8'h00;
            15'd6299: data <= 8'h00;
            15'd6300: data <= 8'h00;
            15'd6301: data <= 8'h00;
            15'd6302: data <= 8'h00;
            15'd6303: data <= 8'h00;
            15'd6304: data <= 8'h01;
            15'd6305: data <= 8'hFF;
            15'd6306: data <= 8'hFF;
            15'd6307: data <= 8'hFF;
            15'd6308: data <= 8'hFF;
            15'd6309: data <= 8'hFF;
            15'd6310: data <= 8'hFF;
            15'd6311: data <= 8'hFF;
            15'd6312: data <= 8'hFF;
            15'd6313: data <= 8'hFF;
            15'd6314: data <= 8'hFF;
            15'd6315: data <= 8'hFF;
            15'd6316: data <= 8'hFF;
            15'd6317: data <= 8'hFF;
            15'd6318: data <= 8'hFF;
            15'd6319: data <= 8'hFF;
            15'd6320: data <= 8'hFF;
            15'd6321: data <= 8'hFF;
            15'd6322: data <= 8'hFF;
            15'd6323: data <= 8'hFF;
            15'd6324: data <= 8'hFF;
            15'd6325: data <= 8'h80;
            15'd6326: data <= 8'h00;
            15'd6327: data <= 8'h00;
            15'd6328: data <= 8'h00;
            15'd6329: data <= 8'h00;
            15'd6330: data <= 8'h00;
            15'd6331: data <= 8'h00;
            15'd6332: data <= 8'h00;
            15'd6333: data <= 8'h00;
            15'd6334: data <= 8'h01;
            15'd6335: data <= 8'hFF;
            15'd6336: data <= 8'hFF;
            15'd6337: data <= 8'hFF;
            15'd6338: data <= 8'hFF;
            15'd6339: data <= 8'hFF;
            15'd6340: data <= 8'hFF;
            15'd6341: data <= 8'hFF;
            15'd6342: data <= 8'hFF;
            15'd6343: data <= 8'hFF;
            15'd6344: data <= 8'hFF;
            15'd6345: data <= 8'hFF;
            15'd6346: data <= 8'hFF;
            15'd6347: data <= 8'hFF;
            15'd6348: data <= 8'hFF;
            15'd6349: data <= 8'hFF;
            15'd6350: data <= 8'hFF;
            15'd6351: data <= 8'hFF;
            15'd6352: data <= 8'hFF;
            15'd6353: data <= 8'hFF;
            15'd6354: data <= 8'hFF;
            15'd6355: data <= 8'h80;
            15'd6356: data <= 8'h00;
            15'd6357: data <= 8'h00;
            15'd6358: data <= 8'h00;
            15'd6359: data <= 8'h00;
            15'd6360: data <= 8'h00;
            15'd6361: data <= 8'h00;
            15'd6362: data <= 8'h00;
            15'd6363: data <= 8'h00;
            15'd6364: data <= 8'h01;
            15'd6365: data <= 8'hFF;
            15'd6366: data <= 8'hFF;
            15'd6367: data <= 8'hFF;
            15'd6368: data <= 8'hFF;
            15'd6369: data <= 8'hFF;
            15'd6370: data <= 8'hFF;
            15'd6371: data <= 8'hFF;
            15'd6372: data <= 8'hFF;
            15'd6373: data <= 8'hFF;
            15'd6374: data <= 8'hFF;
            15'd6375: data <= 8'hFF;
            15'd6376: data <= 8'hFF;
            15'd6377: data <= 8'hFF;
            15'd6378: data <= 8'hFF;
            15'd6379: data <= 8'hFF;
            15'd6380: data <= 8'hFF;
            15'd6381: data <= 8'hFF;
            15'd6382: data <= 8'hFF;
            15'd6383: data <= 8'hFF;
            15'd6384: data <= 8'hFF;
            15'd6385: data <= 8'h80;
            15'd6386: data <= 8'h00;
            15'd6387: data <= 8'h00;
            15'd6388: data <= 8'h00;
            15'd6389: data <= 8'h00;
            15'd6390: data <= 8'h00;
            15'd6391: data <= 8'h00;
            15'd6392: data <= 8'h00;
            15'd6393: data <= 8'h00;
            15'd6394: data <= 8'h01;
            15'd6395: data <= 8'hFF;
            15'd6396: data <= 8'hFF;
            15'd6397: data <= 8'hFF;
            15'd6398: data <= 8'hFF;
            15'd6399: data <= 8'hFF;
            15'd6400: data <= 8'hFF;
            15'd6401: data <= 8'hFF;
            15'd6402: data <= 8'hFF;
            15'd6403: data <= 8'hFF;
            15'd6404: data <= 8'hFF;
            15'd6405: data <= 8'hFF;
            15'd6406: data <= 8'hFF;
            15'd6407: data <= 8'hFF;
            15'd6408: data <= 8'hFF;
            15'd6409: data <= 8'hFF;
            15'd6410: data <= 8'hFF;
            15'd6411: data <= 8'hFF;
            15'd6412: data <= 8'hFF;
            15'd6413: data <= 8'hFF;
            15'd6414: data <= 8'hFF;
            15'd6415: data <= 8'h80;
            15'd6416: data <= 8'h00;
            15'd6417: data <= 8'h00;
            15'd6418: data <= 8'h00;
            15'd6419: data <= 8'h00;
            15'd6420: data <= 8'h00;
            15'd6421: data <= 8'h00;
            15'd6422: data <= 8'h00;
            15'd6423: data <= 8'h00;
            15'd6424: data <= 8'h01;
            15'd6425: data <= 8'hFF;
            15'd6426: data <= 8'hFF;
            15'd6427: data <= 8'hFF;
            15'd6428: data <= 8'hFF;
            15'd6429: data <= 8'hFF;
            15'd6430: data <= 8'hFF;
            15'd6431: data <= 8'hFF;
            15'd6432: data <= 8'hFF;
            15'd6433: data <= 8'hFF;
            15'd6434: data <= 8'hFF;
            15'd6435: data <= 8'hFF;
            15'd6436: data <= 8'hFF;
            15'd6437: data <= 8'hFF;
            15'd6438: data <= 8'hFF;
            15'd6439: data <= 8'hFF;
            15'd6440: data <= 8'hFF;
            15'd6441: data <= 8'hFF;
            15'd6442: data <= 8'hFF;
            15'd6443: data <= 8'hFF;
            15'd6444: data <= 8'hFF;
            15'd6445: data <= 8'h80;
            15'd6446: data <= 8'h00;
            15'd6447: data <= 8'h00;
            15'd6448: data <= 8'h00;
            15'd6449: data <= 8'h00;
            15'd6450: data <= 8'h00;
            15'd6451: data <= 8'h00;
            15'd6452: data <= 8'h00;
            15'd6453: data <= 8'h00;
            15'd6454: data <= 8'h01;
            15'd6455: data <= 8'hFF;
            15'd6456: data <= 8'hFF;
            15'd6457: data <= 8'hFF;
            15'd6458: data <= 8'hFF;
            15'd6459: data <= 8'hFF;
            15'd6460: data <= 8'hFF;
            15'd6461: data <= 8'hFF;
            15'd6462: data <= 8'hFF;
            15'd6463: data <= 8'hFF;
            15'd6464: data <= 8'hFF;
            15'd6465: data <= 8'hFF;
            15'd6466: data <= 8'hFF;
            15'd6467: data <= 8'hFF;
            15'd6468: data <= 8'hFF;
            15'd6469: data <= 8'hFF;
            15'd6470: data <= 8'hFF;
            15'd6471: data <= 8'hFF;
            15'd6472: data <= 8'hFF;
            15'd6473: data <= 8'hFF;
            15'd6474: data <= 8'hFF;
            15'd6475: data <= 8'h80;
            15'd6476: data <= 8'h00;
            15'd6477: data <= 8'h00;
            15'd6478: data <= 8'h00;
            15'd6479: data <= 8'h00;
            15'd6480: data <= 8'h00;
            15'd6481: data <= 8'h00;
            15'd6482: data <= 8'h00;
            15'd6483: data <= 8'h00;
            15'd6484: data <= 8'h01;
            15'd6485: data <= 8'hFF;
            15'd6486: data <= 8'hFF;
            15'd6487: data <= 8'hFF;
            15'd6488: data <= 8'hFF;
            15'd6489: data <= 8'hFF;
            15'd6490: data <= 8'hFF;
            15'd6491: data <= 8'hFF;
            15'd6492: data <= 8'hFF;
            15'd6493: data <= 8'hFF;
            15'd6494: data <= 8'hFF;
            15'd6495: data <= 8'hFF;
            15'd6496: data <= 8'hFF;
            15'd6497: data <= 8'hFF;
            15'd6498: data <= 8'hFF;
            15'd6499: data <= 8'hFF;
            15'd6500: data <= 8'hFF;
            15'd6501: data <= 8'hFF;
            15'd6502: data <= 8'hFF;
            15'd6503: data <= 8'hFF;
            15'd6504: data <= 8'hFF;
            15'd6505: data <= 8'h80;
            15'd6506: data <= 8'h00;
            15'd6507: data <= 8'h00;
            15'd6508: data <= 8'h00;
            15'd6509: data <= 8'h00;
            15'd6510: data <= 8'h00;
            15'd6511: data <= 8'h00;
            15'd6512: data <= 8'h00;
            15'd6513: data <= 8'h00;
            15'd6514: data <= 8'h01;
            15'd6515: data <= 8'hFF;
            15'd6516: data <= 8'hFF;
            15'd6517: data <= 8'hFF;
            15'd6518: data <= 8'hFF;
            15'd6519: data <= 8'hFF;
            15'd6520: data <= 8'hFF;
            15'd6521: data <= 8'hFF;
            15'd6522: data <= 8'hFF;
            15'd6523: data <= 8'hFF;
            15'd6524: data <= 8'hFF;
            15'd6525: data <= 8'hFF;
            15'd6526: data <= 8'hFF;
            15'd6527: data <= 8'hFF;
            15'd6528: data <= 8'hFF;
            15'd6529: data <= 8'hFF;
            15'd6530: data <= 8'hFF;
            15'd6531: data <= 8'hFF;
            15'd6532: data <= 8'hFF;
            15'd6533: data <= 8'hFF;
            15'd6534: data <= 8'hFF;
            15'd6535: data <= 8'h80;
            15'd6536: data <= 8'h00;
            15'd6537: data <= 8'h00;
            15'd6538: data <= 8'h00;
            15'd6539: data <= 8'h00;
            15'd6540: data <= 8'h00;
            15'd6541: data <= 8'h00;
            15'd6542: data <= 8'h00;
            15'd6543: data <= 8'h00;
            15'd6544: data <= 8'h01;
            15'd6545: data <= 8'hFF;
            15'd6546: data <= 8'hFF;
            15'd6547: data <= 8'hFF;
            15'd6548: data <= 8'hFF;
            15'd6549: data <= 8'hFF;
            15'd6550: data <= 8'hFF;
            15'd6551: data <= 8'hFF;
            15'd6552: data <= 8'hFF;
            15'd6553: data <= 8'hFF;
            15'd6554: data <= 8'hFF;
            15'd6555: data <= 8'hFF;
            15'd6556: data <= 8'hFF;
            15'd6557: data <= 8'hFF;
            15'd6558: data <= 8'hFF;
            15'd6559: data <= 8'hFF;
            15'd6560: data <= 8'hFF;
            15'd6561: data <= 8'hFF;
            15'd6562: data <= 8'hFF;
            15'd6563: data <= 8'hFF;
            15'd6564: data <= 8'hFF;
            15'd6565: data <= 8'h80;
            15'd6566: data <= 8'h00;
            15'd6567: data <= 8'h00;
            15'd6568: data <= 8'h00;
            15'd6569: data <= 8'h00;
            15'd6570: data <= 8'h00;
            15'd6571: data <= 8'h00;
            15'd6572: data <= 8'h00;
            15'd6573: data <= 8'h00;
            15'd6574: data <= 8'h01;
            15'd6575: data <= 8'hFF;
            15'd6576: data <= 8'hFF;
            15'd6577: data <= 8'hFF;
            15'd6578: data <= 8'hFF;
            15'd6579: data <= 8'hFF;
            15'd6580: data <= 8'hFF;
            15'd6581: data <= 8'hFF;
            15'd6582: data <= 8'hFF;
            15'd6583: data <= 8'hFF;
            15'd6584: data <= 8'hFF;
            15'd6585: data <= 8'hFF;
            15'd6586: data <= 8'hFF;
            15'd6587: data <= 8'hFF;
            15'd6588: data <= 8'hFF;
            15'd6589: data <= 8'hFF;
            15'd6590: data <= 8'hFF;
            15'd6591: data <= 8'hFF;
            15'd6592: data <= 8'hFF;
            15'd6593: data <= 8'hFF;
            15'd6594: data <= 8'hFF;
            15'd6595: data <= 8'h80;
            15'd6596: data <= 8'h00;
            15'd6597: data <= 8'h00;
            15'd6598: data <= 8'h00;
            15'd6599: data <= 8'h00;
            15'd6600: data <= 8'h00;
            15'd6601: data <= 8'h00;
            15'd6602: data <= 8'h00;
            15'd6603: data <= 8'h00;
            15'd6604: data <= 8'h01;
            15'd6605: data <= 8'hFF;
            15'd6606: data <= 8'hFF;
            15'd6607: data <= 8'hFF;
            15'd6608: data <= 8'hFF;
            15'd6609: data <= 8'hFF;
            15'd6610: data <= 8'hFF;
            15'd6611: data <= 8'hFF;
            15'd6612: data <= 8'hFF;
            15'd6613: data <= 8'hFF;
            15'd6614: data <= 8'hFF;
            15'd6615: data <= 8'hFF;
            15'd6616: data <= 8'hFF;
            15'd6617: data <= 8'hFF;
            15'd6618: data <= 8'hFF;
            15'd6619: data <= 8'hFF;
            15'd6620: data <= 8'hFF;
            15'd6621: data <= 8'hFF;
            15'd6622: data <= 8'hFF;
            15'd6623: data <= 8'hFF;
            15'd6624: data <= 8'hFF;
            15'd6625: data <= 8'h80;
            15'd6626: data <= 8'h00;
            15'd6627: data <= 8'h00;
            15'd6628: data <= 8'h00;
            15'd6629: data <= 8'h00;
            15'd6630: data <= 8'h00;
            15'd6631: data <= 8'h00;
            15'd6632: data <= 8'h00;
            15'd6633: data <= 8'h00;
            15'd6634: data <= 8'h01;
            15'd6635: data <= 8'hFF;
            15'd6636: data <= 8'hFF;
            15'd6637: data <= 8'hFF;
            15'd6638: data <= 8'hFF;
            15'd6639: data <= 8'hFF;
            15'd6640: data <= 8'hFF;
            15'd6641: data <= 8'hFF;
            15'd6642: data <= 8'hFF;
            15'd6643: data <= 8'hFF;
            15'd6644: data <= 8'hFF;
            15'd6645: data <= 8'hFF;
            15'd6646: data <= 8'hFF;
            15'd6647: data <= 8'hFF;
            15'd6648: data <= 8'hFF;
            15'd6649: data <= 8'hFF;
            15'd6650: data <= 8'hFF;
            15'd6651: data <= 8'hFF;
            15'd6652: data <= 8'hFF;
            15'd6653: data <= 8'hFF;
            15'd6654: data <= 8'hFF;
            15'd6655: data <= 8'h80;
            15'd6656: data <= 8'h00;
            15'd6657: data <= 8'h00;
            15'd6658: data <= 8'h00;
            15'd6659: data <= 8'h00;
            15'd6660: data <= 8'h00;
            15'd6661: data <= 8'h00;
            15'd6662: data <= 8'h00;
            15'd6663: data <= 8'h00;
            15'd6664: data <= 8'h01;
            15'd6665: data <= 8'hFF;
            15'd6666: data <= 8'hFF;
            15'd6667: data <= 8'hFF;
            15'd6668: data <= 8'hFF;
            15'd6669: data <= 8'hFF;
            15'd6670: data <= 8'hFF;
            15'd6671: data <= 8'hFF;
            15'd6672: data <= 8'hFF;
            15'd6673: data <= 8'hFF;
            15'd6674: data <= 8'hFF;
            15'd6675: data <= 8'hFF;
            15'd6676: data <= 8'hFF;
            15'd6677: data <= 8'hFF;
            15'd6678: data <= 8'hFF;
            15'd6679: data <= 8'hFF;
            15'd6680: data <= 8'hFF;
            15'd6681: data <= 8'hFF;
            15'd6682: data <= 8'hFF;
            15'd6683: data <= 8'hFF;
            15'd6684: data <= 8'hFF;
            15'd6685: data <= 8'h80;
            15'd6686: data <= 8'h00;
            15'd6687: data <= 8'h00;
            15'd6688: data <= 8'h00;
            15'd6689: data <= 8'h00;
            15'd6690: data <= 8'h00;
            15'd6691: data <= 8'h00;
            15'd6692: data <= 8'h00;
            15'd6693: data <= 8'h00;
            15'd6694: data <= 8'h01;
            15'd6695: data <= 8'hFF;
            15'd6696: data <= 8'hFF;
            15'd6697: data <= 8'hFF;
            15'd6698: data <= 8'hFF;
            15'd6699: data <= 8'hFF;
            15'd6700: data <= 8'hFF;
            15'd6701: data <= 8'hFF;
            15'd6702: data <= 8'hFF;
            15'd6703: data <= 8'hFF;
            15'd6704: data <= 8'hFF;
            15'd6705: data <= 8'hFF;
            15'd6706: data <= 8'hFF;
            15'd6707: data <= 8'hFF;
            15'd6708: data <= 8'hFF;
            15'd6709: data <= 8'hFF;
            15'd6710: data <= 8'hFF;
            15'd6711: data <= 8'hFF;
            15'd6712: data <= 8'hFF;
            15'd6713: data <= 8'hFF;
            15'd6714: data <= 8'hFF;
            15'd6715: data <= 8'h80;
            15'd6716: data <= 8'h00;
            15'd6717: data <= 8'h00;
            15'd6718: data <= 8'h00;
            15'd6719: data <= 8'h00;
            15'd6720: data <= 8'h00;
            15'd6721: data <= 8'h00;
            15'd6722: data <= 8'h00;
            15'd6723: data <= 8'h00;
            15'd6724: data <= 8'h01;
            15'd6725: data <= 8'hFF;
            15'd6726: data <= 8'hFF;
            15'd6727: data <= 8'hFF;
            15'd6728: data <= 8'hFF;
            15'd6729: data <= 8'hFF;
            15'd6730: data <= 8'hFF;
            15'd6731: data <= 8'hFF;
            15'd6732: data <= 8'hFF;
            15'd6733: data <= 8'hFF;
            15'd6734: data <= 8'hFF;
            15'd6735: data <= 8'hFF;
            15'd6736: data <= 8'hFF;
            15'd6737: data <= 8'hFF;
            15'd6738: data <= 8'hFF;
            15'd6739: data <= 8'hFF;
            15'd6740: data <= 8'hFF;
            15'd6741: data <= 8'hFF;
            15'd6742: data <= 8'hFF;
            15'd6743: data <= 8'hFF;
            15'd6744: data <= 8'hFF;
            15'd6745: data <= 8'h80;
            15'd6746: data <= 8'h00;
            15'd6747: data <= 8'h00;
            15'd6748: data <= 8'h00;
            15'd6749: data <= 8'h00;
            15'd6750: data <= 8'h00;
            15'd6751: data <= 8'h00;
            15'd6752: data <= 8'h00;
            15'd6753: data <= 8'h00;
            15'd6754: data <= 8'h01;
            15'd6755: data <= 8'hFF;
            15'd6756: data <= 8'hFF;
            15'd6757: data <= 8'hFF;
            15'd6758: data <= 8'hFF;
            15'd6759: data <= 8'hFF;
            15'd6760: data <= 8'hFF;
            15'd6761: data <= 8'hFF;
            15'd6762: data <= 8'hFF;
            15'd6763: data <= 8'hFF;
            15'd6764: data <= 8'hFF;
            15'd6765: data <= 8'hFF;
            15'd6766: data <= 8'hFF;
            15'd6767: data <= 8'hFF;
            15'd6768: data <= 8'hFF;
            15'd6769: data <= 8'hFF;
            15'd6770: data <= 8'hFF;
            15'd6771: data <= 8'hFF;
            15'd6772: data <= 8'hFF;
            15'd6773: data <= 8'hFF;
            15'd6774: data <= 8'hFF;
            15'd6775: data <= 8'h80;
            15'd6776: data <= 8'h00;
            15'd6777: data <= 8'h00;
            15'd6778: data <= 8'h00;
            15'd6779: data <= 8'h00;
            15'd6780: data <= 8'h00;
            15'd6781: data <= 8'h00;
            15'd6782: data <= 8'h00;
            15'd6783: data <= 8'h00;
            15'd6784: data <= 8'h01;
            15'd6785: data <= 8'hFF;
            15'd6786: data <= 8'hFF;
            15'd6787: data <= 8'hFF;
            15'd6788: data <= 8'hFF;
            15'd6789: data <= 8'hFF;
            15'd6790: data <= 8'hFF;
            15'd6791: data <= 8'hFF;
            15'd6792: data <= 8'hFF;
            15'd6793: data <= 8'hFF;
            15'd6794: data <= 8'hFF;
            15'd6795: data <= 8'hFF;
            15'd6796: data <= 8'hFF;
            15'd6797: data <= 8'hF7;
            15'd6798: data <= 8'hFF;
            15'd6799: data <= 8'hFF;
            15'd6800: data <= 8'hFF;
            15'd6801: data <= 8'hFF;
            15'd6802: data <= 8'hFF;
            15'd6803: data <= 8'hFF;
            15'd6804: data <= 8'hFF;
            15'd6805: data <= 8'h80;
            15'd6806: data <= 8'h00;
            15'd6807: data <= 8'h00;
            15'd6808: data <= 8'h00;
            15'd6809: data <= 8'h00;
            15'd6810: data <= 8'h00;
            15'd6811: data <= 8'h00;
            15'd6812: data <= 8'h00;
            15'd6813: data <= 8'h00;
            15'd6814: data <= 8'h01;
            15'd6815: data <= 8'hFF;
            15'd6816: data <= 8'hFF;
            15'd6817: data <= 8'hFF;
            15'd6818: data <= 8'hFF;
            15'd6819: data <= 8'hFF;
            15'd6820: data <= 8'hFF;
            15'd6821: data <= 8'hFF;
            15'd6822: data <= 8'h83;
            15'd6823: data <= 8'hFF;
            15'd6824: data <= 8'hFF;
            15'd6825: data <= 8'hFF;
            15'd6826: data <= 8'hFF;
            15'd6827: data <= 8'h03;
            15'd6828: data <= 8'hFF;
            15'd6829: data <= 8'hFF;
            15'd6830: data <= 8'hFF;
            15'd6831: data <= 8'hFF;
            15'd6832: data <= 8'hFF;
            15'd6833: data <= 8'hFF;
            15'd6834: data <= 8'hFF;
            15'd6835: data <= 8'h80;
            15'd6836: data <= 8'h00;
            15'd6837: data <= 8'h00;
            15'd6838: data <= 8'h00;
            15'd6839: data <= 8'h00;
            15'd6840: data <= 8'h00;
            15'd6841: data <= 8'h00;
            15'd6842: data <= 8'h00;
            15'd6843: data <= 8'h00;
            15'd6844: data <= 8'h01;
            15'd6845: data <= 8'hFF;
            15'd6846: data <= 8'hFF;
            15'd6847: data <= 8'hFF;
            15'd6848: data <= 8'hFF;
            15'd6849: data <= 8'hFF;
            15'd6850: data <= 8'hFF;
            15'd6851: data <= 8'hFF;
            15'd6852: data <= 8'h80;
            15'd6853: data <= 8'h7F;
            15'd6854: data <= 8'hFF;
            15'd6855: data <= 8'hFF;
            15'd6856: data <= 8'hFC;
            15'd6857: data <= 8'h03;
            15'd6858: data <= 8'hFF;
            15'd6859: data <= 8'hFF;
            15'd6860: data <= 8'hFF;
            15'd6861: data <= 8'hFF;
            15'd6862: data <= 8'hFF;
            15'd6863: data <= 8'hFF;
            15'd6864: data <= 8'hFF;
            15'd6865: data <= 8'h80;
            15'd6866: data <= 8'h00;
            15'd6867: data <= 8'h00;
            15'd6868: data <= 8'h00;
            15'd6869: data <= 8'h00;
            15'd6870: data <= 8'h00;
            15'd6871: data <= 8'h00;
            15'd6872: data <= 8'h00;
            15'd6873: data <= 8'h00;
            15'd6874: data <= 8'h01;
            15'd6875: data <= 8'hFF;
            15'd6876: data <= 8'hFF;
            15'd6877: data <= 8'hFF;
            15'd6878: data <= 8'hFF;
            15'd6879: data <= 8'hFF;
            15'd6880: data <= 8'hFF;
            15'd6881: data <= 8'hFF;
            15'd6882: data <= 8'h00;
            15'd6883: data <= 8'h07;
            15'd6884: data <= 8'hFF;
            15'd6885: data <= 8'hFF;
            15'd6886: data <= 8'hF8;
            15'd6887: data <= 8'h03;
            15'd6888: data <= 8'hFF;
            15'd6889: data <= 8'hFF;
            15'd6890: data <= 8'hFF;
            15'd6891: data <= 8'hFF;
            15'd6892: data <= 8'hFF;
            15'd6893: data <= 8'hFF;
            15'd6894: data <= 8'hFF;
            15'd6895: data <= 8'h80;
            15'd6896: data <= 8'h00;
            15'd6897: data <= 8'h00;
            15'd6898: data <= 8'h00;
            15'd6899: data <= 8'h00;
            15'd6900: data <= 8'h00;
            15'd6901: data <= 8'h00;
            15'd6902: data <= 8'h00;
            15'd6903: data <= 8'h00;
            15'd6904: data <= 8'h01;
            15'd6905: data <= 8'hFF;
            15'd6906: data <= 8'hFF;
            15'd6907: data <= 8'hFF;
            15'd6908: data <= 8'hFF;
            15'd6909: data <= 8'hFF;
            15'd6910: data <= 8'hFF;
            15'd6911: data <= 8'hFF;
            15'd6912: data <= 8'h80;
            15'd6913: data <= 8'h01;
            15'd6914: data <= 8'hFF;
            15'd6915: data <= 8'hFF;
            15'd6916: data <= 8'hE0;
            15'd6917: data <= 8'h07;
            15'd6918: data <= 8'hFF;
            15'd6919: data <= 8'hFF;
            15'd6920: data <= 8'hFF;
            15'd6921: data <= 8'hFF;
            15'd6922: data <= 8'hFF;
            15'd6923: data <= 8'hFF;
            15'd6924: data <= 8'hFF;
            15'd6925: data <= 8'h80;
            15'd6926: data <= 8'h00;
            15'd6927: data <= 8'h00;
            15'd6928: data <= 8'h00;
            15'd6929: data <= 8'h00;
            15'd6930: data <= 8'h00;
            15'd6931: data <= 8'h00;
            15'd6932: data <= 8'h00;
            15'd6933: data <= 8'h00;
            15'd6934: data <= 8'h01;
            15'd6935: data <= 8'hFF;
            15'd6936: data <= 8'hFF;
            15'd6937: data <= 8'hFF;
            15'd6938: data <= 8'hFF;
            15'd6939: data <= 8'hFF;
            15'd6940: data <= 8'hFF;
            15'd6941: data <= 8'hFF;
            15'd6942: data <= 8'hE0;
            15'd6943: data <= 8'h00;
            15'd6944: data <= 8'hFF;
            15'd6945: data <= 8'hFF;
            15'd6946: data <= 8'hC0;
            15'd6947: data <= 8'h1F;
            15'd6948: data <= 8'hFF;
            15'd6949: data <= 8'hFF;
            15'd6950: data <= 8'hFF;
            15'd6951: data <= 8'hFF;
            15'd6952: data <= 8'hFF;
            15'd6953: data <= 8'hFF;
            15'd6954: data <= 8'hFF;
            15'd6955: data <= 8'h80;
            15'd6956: data <= 8'h00;
            15'd6957: data <= 8'h00;
            15'd6958: data <= 8'h00;
            15'd6959: data <= 8'h00;
            15'd6960: data <= 8'h00;
            15'd6961: data <= 8'h00;
            15'd6962: data <= 8'h00;
            15'd6963: data <= 8'h00;
            15'd6964: data <= 8'h01;
            15'd6965: data <= 8'hFF;
            15'd6966: data <= 8'hFF;
            15'd6967: data <= 8'hFF;
            15'd6968: data <= 8'hFF;
            15'd6969: data <= 8'hFF;
            15'd6970: data <= 8'hFF;
            15'd6971: data <= 8'hFF;
            15'd6972: data <= 8'hFC;
            15'd6973: data <= 8'h00;
            15'd6974: data <= 8'h7F;
            15'd6975: data <= 8'hFF;
            15'd6976: data <= 8'h00;
            15'd6977: data <= 8'h7F;
            15'd6978: data <= 8'hFF;
            15'd6979: data <= 8'hFF;
            15'd6980: data <= 8'hFF;
            15'd6981: data <= 8'hFF;
            15'd6982: data <= 8'hFF;
            15'd6983: data <= 8'hFF;
            15'd6984: data <= 8'hFF;
            15'd6985: data <= 8'h80;
            15'd6986: data <= 8'h00;
            15'd6987: data <= 8'h00;
            15'd6988: data <= 8'h00;
            15'd6989: data <= 8'h00;
            15'd6990: data <= 8'h00;
            15'd6991: data <= 8'h00;
            15'd6992: data <= 8'h00;
            15'd6993: data <= 8'h00;
            15'd6994: data <= 8'h01;
            15'd6995: data <= 8'hFF;
            15'd6996: data <= 8'hFF;
            15'd6997: data <= 8'hFF;
            15'd6998: data <= 8'hFF;
            15'd6999: data <= 8'hFF;
            15'd7000: data <= 8'hFF;
            15'd7001: data <= 8'hFF;
            15'd7002: data <= 8'hFF;
            15'd7003: data <= 8'h00;
            15'd7004: data <= 8'hFF;
            15'd7005: data <= 8'hFF;
            15'd7006: data <= 8'h01;
            15'd7007: data <= 8'hFF;
            15'd7008: data <= 8'hFF;
            15'd7009: data <= 8'hFF;
            15'd7010: data <= 8'hFF;
            15'd7011: data <= 8'hFF;
            15'd7012: data <= 8'hFF;
            15'd7013: data <= 8'hFF;
            15'd7014: data <= 8'hFF;
            15'd7015: data <= 8'h80;
            15'd7016: data <= 8'h00;
            15'd7017: data <= 8'h00;
            15'd7018: data <= 8'h00;
            15'd7019: data <= 8'h00;
            15'd7020: data <= 8'h00;
            15'd7021: data <= 8'h00;
            15'd7022: data <= 8'h00;
            15'd7023: data <= 8'h00;
            15'd7024: data <= 8'h01;
            15'd7025: data <= 8'hFF;
            15'd7026: data <= 8'hFF;
            15'd7027: data <= 8'hFF;
            15'd7028: data <= 8'hFF;
            15'd7029: data <= 8'hFF;
            15'd7030: data <= 8'hFF;
            15'd7031: data <= 8'hFF;
            15'd7032: data <= 8'hFF;
            15'd7033: data <= 8'hF1;
            15'd7034: data <= 8'hFF;
            15'd7035: data <= 8'hFE;
            15'd7036: data <= 8'h07;
            15'd7037: data <= 8'hFF;
            15'd7038: data <= 8'hFF;
            15'd7039: data <= 8'hFF;
            15'd7040: data <= 8'hFF;
            15'd7041: data <= 8'hFF;
            15'd7042: data <= 8'hFF;
            15'd7043: data <= 8'hFF;
            15'd7044: data <= 8'hFF;
            15'd7045: data <= 8'h80;
            15'd7046: data <= 8'h00;
            15'd7047: data <= 8'h00;
            15'd7048: data <= 8'h00;
            15'd7049: data <= 8'h00;
            15'd7050: data <= 8'h00;
            15'd7051: data <= 8'h00;
            15'd7052: data <= 8'h00;
            15'd7053: data <= 8'h00;
            15'd7054: data <= 8'h01;
            15'd7055: data <= 8'hFF;
            15'd7056: data <= 8'hFF;
            15'd7057: data <= 8'hFF;
            15'd7058: data <= 8'hFF;
            15'd7059: data <= 8'hFF;
            15'd7060: data <= 8'hFF;
            15'd7061: data <= 8'hFF;
            15'd7062: data <= 8'hFF;
            15'd7063: data <= 8'hFF;
            15'd7064: data <= 8'hFF;
            15'd7065: data <= 8'hFF;
            15'd7066: data <= 8'h1F;
            15'd7067: data <= 8'hFF;
            15'd7068: data <= 8'hFF;
            15'd7069: data <= 8'hFF;
            15'd7070: data <= 8'hFF;
            15'd7071: data <= 8'hFF;
            15'd7072: data <= 8'hFF;
            15'd7073: data <= 8'hFF;
            15'd7074: data <= 8'hFF;
            15'd7075: data <= 8'h80;
            15'd7076: data <= 8'h00;
            15'd7077: data <= 8'h00;
            15'd7078: data <= 8'h00;
            15'd7079: data <= 8'h00;
            15'd7080: data <= 8'h00;
            15'd7081: data <= 8'h00;
            15'd7082: data <= 8'h00;
            15'd7083: data <= 8'h00;
            15'd7084: data <= 8'h01;
            15'd7085: data <= 8'hFF;
            15'd7086: data <= 8'hFF;
            15'd7087: data <= 8'hFF;
            15'd7088: data <= 8'hFF;
            15'd7089: data <= 8'hFF;
            15'd7090: data <= 8'hFF;
            15'd7091: data <= 8'hFF;
            15'd7092: data <= 8'hFF;
            15'd7093: data <= 8'hFF;
            15'd7094: data <= 8'hFF;
            15'd7095: data <= 8'hFF;
            15'd7096: data <= 8'hFF;
            15'd7097: data <= 8'hFF;
            15'd7098: data <= 8'hFF;
            15'd7099: data <= 8'hFF;
            15'd7100: data <= 8'hFF;
            15'd7101: data <= 8'hFF;
            15'd7102: data <= 8'hFF;
            15'd7103: data <= 8'hFF;
            15'd7104: data <= 8'hFF;
            15'd7105: data <= 8'h80;
            15'd7106: data <= 8'h00;
            15'd7107: data <= 8'h00;
            15'd7108: data <= 8'h00;
            15'd7109: data <= 8'h00;
            15'd7110: data <= 8'h00;
            15'd7111: data <= 8'h00;
            15'd7112: data <= 8'h00;
            15'd7113: data <= 8'h00;
            15'd7114: data <= 8'h01;
            15'd7115: data <= 8'hFF;
            15'd7116: data <= 8'hFF;
            15'd7117: data <= 8'hFF;
            15'd7118: data <= 8'hFF;
            15'd7119: data <= 8'hFF;
            15'd7120: data <= 8'hFF;
            15'd7121: data <= 8'hFF;
            15'd7122: data <= 8'hFF;
            15'd7123: data <= 8'hFF;
            15'd7124: data <= 8'hFF;
            15'd7125: data <= 8'hFF;
            15'd7126: data <= 8'hFF;
            15'd7127: data <= 8'hFF;
            15'd7128: data <= 8'hFF;
            15'd7129: data <= 8'hFF;
            15'd7130: data <= 8'hFF;
            15'd7131: data <= 8'hFF;
            15'd7132: data <= 8'hFF;
            15'd7133: data <= 8'hFF;
            15'd7134: data <= 8'hFF;
            15'd7135: data <= 8'h80;
            15'd7136: data <= 8'h00;
            15'd7137: data <= 8'h00;
            15'd7138: data <= 8'h00;
            15'd7139: data <= 8'h00;
            15'd7140: data <= 8'h00;
            15'd7141: data <= 8'h00;
            15'd7142: data <= 8'h00;
            15'd7143: data <= 8'h00;
            15'd7144: data <= 8'h01;
            15'd7145: data <= 8'hFF;
            15'd7146: data <= 8'hFF;
            15'd7147: data <= 8'hFF;
            15'd7148: data <= 8'hFF;
            15'd7149: data <= 8'hFF;
            15'd7150: data <= 8'hFF;
            15'd7151: data <= 8'hFF;
            15'd7152: data <= 8'hFF;
            15'd7153: data <= 8'hDF;
            15'd7154: data <= 8'hFF;
            15'd7155: data <= 8'hFF;
            15'd7156: data <= 8'hFF;
            15'd7157: data <= 8'hFF;
            15'd7158: data <= 8'hFF;
            15'd7159: data <= 8'hFF;
            15'd7160: data <= 8'hFF;
            15'd7161: data <= 8'hFF;
            15'd7162: data <= 8'hFF;
            15'd7163: data <= 8'hFF;
            15'd7164: data <= 8'hFF;
            15'd7165: data <= 8'h80;
            15'd7166: data <= 8'h00;
            15'd7167: data <= 8'h00;
            15'd7168: data <= 8'h00;
            15'd7169: data <= 8'h00;
            15'd7170: data <= 8'h00;
            15'd7171: data <= 8'h00;
            15'd7172: data <= 8'h00;
            15'd7173: data <= 8'h00;
            15'd7174: data <= 8'h01;
            15'd7175: data <= 8'hFF;
            15'd7176: data <= 8'hFF;
            15'd7177: data <= 8'hFF;
            15'd7178: data <= 8'hFF;
            15'd7179: data <= 8'hFF;
            15'd7180: data <= 8'hFF;
            15'd7181: data <= 8'hFF;
            15'd7182: data <= 8'hFF;
            15'd7183: data <= 8'h07;
            15'd7184: data <= 8'hFF;
            15'd7185: data <= 8'hFF;
            15'd7186: data <= 8'hF0;
            15'd7187: data <= 8'h7F;
            15'd7188: data <= 8'hFF;
            15'd7189: data <= 8'hFF;
            15'd7190: data <= 8'hFF;
            15'd7191: data <= 8'hFF;
            15'd7192: data <= 8'hFF;
            15'd7193: data <= 8'hFF;
            15'd7194: data <= 8'hFF;
            15'd7195: data <= 8'h80;
            15'd7196: data <= 8'h00;
            15'd7197: data <= 8'h00;
            15'd7198: data <= 8'h00;
            15'd7199: data <= 8'h00;
            15'd7200: data <= 8'h00;
            15'd7201: data <= 8'h00;
            15'd7202: data <= 8'h00;
            15'd7203: data <= 8'h00;
            15'd7204: data <= 8'h01;
            15'd7205: data <= 8'hFF;
            15'd7206: data <= 8'hFF;
            15'd7207: data <= 8'hFF;
            15'd7208: data <= 8'hFF;
            15'd7209: data <= 8'hFF;
            15'd7210: data <= 8'hFF;
            15'd7211: data <= 8'hFF;
            15'd7212: data <= 8'hFE;
            15'd7213: data <= 8'h07;
            15'd7214: data <= 8'hFF;
            15'd7215: data <= 8'hFF;
            15'd7216: data <= 8'hE0;
            15'd7217: data <= 8'h7F;
            15'd7218: data <= 8'hFF;
            15'd7219: data <= 8'hFF;
            15'd7220: data <= 8'hFF;
            15'd7221: data <= 8'hFF;
            15'd7222: data <= 8'hFF;
            15'd7223: data <= 8'hFF;
            15'd7224: data <= 8'hFF;
            15'd7225: data <= 8'h80;
            15'd7226: data <= 8'h00;
            15'd7227: data <= 8'h00;
            15'd7228: data <= 8'h00;
            15'd7229: data <= 8'h00;
            15'd7230: data <= 8'h00;
            15'd7231: data <= 8'h00;
            15'd7232: data <= 8'h00;
            15'd7233: data <= 8'h00;
            15'd7234: data <= 8'h01;
            15'd7235: data <= 8'hFF;
            15'd7236: data <= 8'hFF;
            15'd7237: data <= 8'hFF;
            15'd7238: data <= 8'hFF;
            15'd7239: data <= 8'hFF;
            15'd7240: data <= 8'hFF;
            15'd7241: data <= 8'hFF;
            15'd7242: data <= 8'hFC;
            15'd7243: data <= 8'h03;
            15'd7244: data <= 8'hFF;
            15'd7245: data <= 8'hFF;
            15'd7246: data <= 8'hC0;
            15'd7247: data <= 8'h3F;
            15'd7248: data <= 8'hFF;
            15'd7249: data <= 8'hFF;
            15'd7250: data <= 8'hFF;
            15'd7251: data <= 8'hFF;
            15'd7252: data <= 8'hFF;
            15'd7253: data <= 8'hFF;
            15'd7254: data <= 8'hFF;
            15'd7255: data <= 8'h80;
            15'd7256: data <= 8'h00;
            15'd7257: data <= 8'h00;
            15'd7258: data <= 8'h00;
            15'd7259: data <= 8'h00;
            15'd7260: data <= 8'h00;
            15'd7261: data <= 8'h00;
            15'd7262: data <= 8'h00;
            15'd7263: data <= 8'h00;
            15'd7264: data <= 8'h01;
            15'd7265: data <= 8'hFF;
            15'd7266: data <= 8'hFF;
            15'd7267: data <= 8'hFF;
            15'd7268: data <= 8'hFF;
            15'd7269: data <= 8'hFF;
            15'd7270: data <= 8'hFF;
            15'd7271: data <= 8'hFF;
            15'd7272: data <= 8'hFC;
            15'd7273: data <= 8'h03;
            15'd7274: data <= 8'hFF;
            15'd7275: data <= 8'hFF;
            15'd7276: data <= 8'hC0;
            15'd7277: data <= 8'h3F;
            15'd7278: data <= 8'hFF;
            15'd7279: data <= 8'hFF;
            15'd7280: data <= 8'hFF;
            15'd7281: data <= 8'hFF;
            15'd7282: data <= 8'hFF;
            15'd7283: data <= 8'hFF;
            15'd7284: data <= 8'hFF;
            15'd7285: data <= 8'h80;
            15'd7286: data <= 8'h00;
            15'd7287: data <= 8'h00;
            15'd7288: data <= 8'h00;
            15'd7289: data <= 8'h00;
            15'd7290: data <= 8'h00;
            15'd7291: data <= 8'h00;
            15'd7292: data <= 8'h00;
            15'd7293: data <= 8'h00;
            15'd7294: data <= 8'h01;
            15'd7295: data <= 8'hFF;
            15'd7296: data <= 8'hFF;
            15'd7297: data <= 8'hFF;
            15'd7298: data <= 8'hFF;
            15'd7299: data <= 8'hFF;
            15'd7300: data <= 8'hFF;
            15'd7301: data <= 8'hFF;
            15'd7302: data <= 8'hFC;
            15'd7303: data <= 8'h03;
            15'd7304: data <= 8'hFF;
            15'd7305: data <= 8'hFF;
            15'd7306: data <= 8'hC0;
            15'd7307: data <= 8'h3F;
            15'd7308: data <= 8'hFF;
            15'd7309: data <= 8'hFF;
            15'd7310: data <= 8'hFF;
            15'd7311: data <= 8'hFF;
            15'd7312: data <= 8'hFF;
            15'd7313: data <= 8'hFF;
            15'd7314: data <= 8'hFF;
            15'd7315: data <= 8'h80;
            15'd7316: data <= 8'h00;
            15'd7317: data <= 8'h00;
            15'd7318: data <= 8'h00;
            15'd7319: data <= 8'h00;
            15'd7320: data <= 8'h00;
            15'd7321: data <= 8'h00;
            15'd7322: data <= 8'h00;
            15'd7323: data <= 8'h00;
            15'd7324: data <= 8'h01;
            15'd7325: data <= 8'hFF;
            15'd7326: data <= 8'hFF;
            15'd7327: data <= 8'hFF;
            15'd7328: data <= 8'hFF;
            15'd7329: data <= 8'hFF;
            15'd7330: data <= 8'hFF;
            15'd7331: data <= 8'hFF;
            15'd7332: data <= 8'hFC;
            15'd7333: data <= 8'h03;
            15'd7334: data <= 8'hFF;
            15'd7335: data <= 8'hFF;
            15'd7336: data <= 8'hC0;
            15'd7337: data <= 8'h7F;
            15'd7338: data <= 8'hFF;
            15'd7339: data <= 8'hFF;
            15'd7340: data <= 8'hFF;
            15'd7341: data <= 8'hFF;
            15'd7342: data <= 8'hFF;
            15'd7343: data <= 8'hFF;
            15'd7344: data <= 8'hFF;
            15'd7345: data <= 8'h80;
            15'd7346: data <= 8'h00;
            15'd7347: data <= 8'h00;
            15'd7348: data <= 8'h00;
            15'd7349: data <= 8'h00;
            15'd7350: data <= 8'h00;
            15'd7351: data <= 8'h00;
            15'd7352: data <= 8'h00;
            15'd7353: data <= 8'h00;
            15'd7354: data <= 8'h01;
            15'd7355: data <= 8'hFF;
            15'd7356: data <= 8'hFF;
            15'd7357: data <= 8'hFF;
            15'd7358: data <= 8'hFF;
            15'd7359: data <= 8'hFF;
            15'd7360: data <= 8'hFF;
            15'd7361: data <= 8'hFF;
            15'd7362: data <= 8'hFE;
            15'd7363: data <= 8'h07;
            15'd7364: data <= 8'hFF;
            15'd7365: data <= 8'hFF;
            15'd7366: data <= 8'hE0;
            15'd7367: data <= 8'h7F;
            15'd7368: data <= 8'hFF;
            15'd7369: data <= 8'hFF;
            15'd7370: data <= 8'hFF;
            15'd7371: data <= 8'hFF;
            15'd7372: data <= 8'hFF;
            15'd7373: data <= 8'hFF;
            15'd7374: data <= 8'hFF;
            15'd7375: data <= 8'h80;
            15'd7376: data <= 8'h00;
            15'd7377: data <= 8'h00;
            15'd7378: data <= 8'h00;
            15'd7379: data <= 8'h00;
            15'd7380: data <= 8'h00;
            15'd7381: data <= 8'h00;
            15'd7382: data <= 8'h00;
            15'd7383: data <= 8'h00;
            15'd7384: data <= 8'h01;
            15'd7385: data <= 8'hFF;
            15'd7386: data <= 8'hFF;
            15'd7387: data <= 8'hFF;
            15'd7388: data <= 8'hFF;
            15'd7389: data <= 8'hFF;
            15'd7390: data <= 8'hFF;
            15'd7391: data <= 8'hFF;
            15'd7392: data <= 8'hFF;
            15'd7393: data <= 8'h1F;
            15'd7394: data <= 8'hFF;
            15'd7395: data <= 8'hFF;
            15'd7396: data <= 8'hF9;
            15'd7397: data <= 8'hFF;
            15'd7398: data <= 8'hFF;
            15'd7399: data <= 8'hFF;
            15'd7400: data <= 8'hFF;
            15'd7401: data <= 8'hFF;
            15'd7402: data <= 8'hFF;
            15'd7403: data <= 8'hFF;
            15'd7404: data <= 8'hFF;
            15'd7405: data <= 8'h80;
            15'd7406: data <= 8'h00;
            15'd7407: data <= 8'h00;
            15'd7408: data <= 8'h00;
            15'd7409: data <= 8'h00;
            15'd7410: data <= 8'h00;
            15'd7411: data <= 8'h00;
            15'd7412: data <= 8'h00;
            15'd7413: data <= 8'h00;
            15'd7414: data <= 8'h01;
            15'd7415: data <= 8'hFF;
            15'd7416: data <= 8'hFF;
            15'd7417: data <= 8'hFF;
            15'd7418: data <= 8'hFF;
            15'd7419: data <= 8'hFF;
            15'd7420: data <= 8'hFF;
            15'd7421: data <= 8'hFF;
            15'd7422: data <= 8'hFF;
            15'd7423: data <= 8'hFF;
            15'd7424: data <= 8'hFF;
            15'd7425: data <= 8'hFF;
            15'd7426: data <= 8'hFF;
            15'd7427: data <= 8'hFF;
            15'd7428: data <= 8'hFF;
            15'd7429: data <= 8'hFF;
            15'd7430: data <= 8'hFF;
            15'd7431: data <= 8'hFF;
            15'd7432: data <= 8'hFF;
            15'd7433: data <= 8'hFF;
            15'd7434: data <= 8'hFF;
            15'd7435: data <= 8'h80;
            15'd7436: data <= 8'h00;
            15'd7437: data <= 8'h00;
            15'd7438: data <= 8'h00;
            15'd7439: data <= 8'h00;
            15'd7440: data <= 8'h00;
            15'd7441: data <= 8'h00;
            15'd7442: data <= 8'h00;
            15'd7443: data <= 8'h00;
            15'd7444: data <= 8'h01;
            15'd7445: data <= 8'hFF;
            15'd7446: data <= 8'hFF;
            15'd7447: data <= 8'hFF;
            15'd7448: data <= 8'hFF;
            15'd7449: data <= 8'hFF;
            15'd7450: data <= 8'hFF;
            15'd7451: data <= 8'hFF;
            15'd7452: data <= 8'hFF;
            15'd7453: data <= 8'hFF;
            15'd7454: data <= 8'hFF;
            15'd7455: data <= 8'hFF;
            15'd7456: data <= 8'hFF;
            15'd7457: data <= 8'hFF;
            15'd7458: data <= 8'hFF;
            15'd7459: data <= 8'hFF;
            15'd7460: data <= 8'hFF;
            15'd7461: data <= 8'hFF;
            15'd7462: data <= 8'hFF;
            15'd7463: data <= 8'hFF;
            15'd7464: data <= 8'hFF;
            15'd7465: data <= 8'h80;
            15'd7466: data <= 8'h00;
            15'd7467: data <= 8'h00;
            15'd7468: data <= 8'h00;
            15'd7469: data <= 8'h00;
            15'd7470: data <= 8'h00;
            15'd7471: data <= 8'h00;
            15'd7472: data <= 8'h00;
            15'd7473: data <= 8'h00;
            15'd7474: data <= 8'h01;
            15'd7475: data <= 8'hFF;
            15'd7476: data <= 8'hFF;
            15'd7477: data <= 8'hFF;
            15'd7478: data <= 8'hFF;
            15'd7479: data <= 8'hFF;
            15'd7480: data <= 8'hFF;
            15'd7481: data <= 8'hFF;
            15'd7482: data <= 8'hFF;
            15'd7483: data <= 8'hFF;
            15'd7484: data <= 8'hFF;
            15'd7485: data <= 8'hFF;
            15'd7486: data <= 8'hFF;
            15'd7487: data <= 8'hFF;
            15'd7488: data <= 8'hFF;
            15'd7489: data <= 8'hFF;
            15'd7490: data <= 8'hFF;
            15'd7491: data <= 8'hFF;
            15'd7492: data <= 8'hFF;
            15'd7493: data <= 8'hFF;
            15'd7494: data <= 8'hFF;
            15'd7495: data <= 8'h80;
            15'd7496: data <= 8'h00;
            15'd7497: data <= 8'h00;
            15'd7498: data <= 8'h00;
            15'd7499: data <= 8'h00;
            15'd7500: data <= 8'h00;
            15'd7501: data <= 8'h00;
            15'd7502: data <= 8'h00;
            15'd7503: data <= 8'h00;
            15'd7504: data <= 8'h01;
            15'd7505: data <= 8'hFF;
            15'd7506: data <= 8'hFF;
            15'd7507: data <= 8'hFF;
            15'd7508: data <= 8'hFF;
            15'd7509: data <= 8'hFF;
            15'd7510: data <= 8'hFF;
            15'd7511: data <= 8'hFF;
            15'd7512: data <= 8'hFF;
            15'd7513: data <= 8'hFF;
            15'd7514: data <= 8'hFF;
            15'd7515: data <= 8'hFF;
            15'd7516: data <= 8'hFF;
            15'd7517: data <= 8'hFF;
            15'd7518: data <= 8'hFF;
            15'd7519: data <= 8'hFF;
            15'd7520: data <= 8'hFF;
            15'd7521: data <= 8'hFF;
            15'd7522: data <= 8'hFF;
            15'd7523: data <= 8'hFF;
            15'd7524: data <= 8'hFF;
            15'd7525: data <= 8'h80;
            15'd7526: data <= 8'h00;
            15'd7527: data <= 8'h00;
            15'd7528: data <= 8'h00;
            15'd7529: data <= 8'h00;
            15'd7530: data <= 8'h00;
            15'd7531: data <= 8'h00;
            15'd7532: data <= 8'h00;
            15'd7533: data <= 8'h00;
            15'd7534: data <= 8'h01;
            15'd7535: data <= 8'hFF;
            15'd7536: data <= 8'hFF;
            15'd7537: data <= 8'hFF;
            15'd7538: data <= 8'hFF;
            15'd7539: data <= 8'hFF;
            15'd7540: data <= 8'hFF;
            15'd7541: data <= 8'hFE;
            15'd7542: data <= 8'h7F;
            15'd7543: data <= 8'hFF;
            15'd7544: data <= 8'hFF;
            15'd7545: data <= 8'hFF;
            15'd7546: data <= 8'hFF;
            15'd7547: data <= 8'hFF;
            15'd7548: data <= 8'hF1;
            15'd7549: data <= 8'hF1;
            15'd7550: data <= 8'hFF;
            15'd7551: data <= 8'hFF;
            15'd7552: data <= 8'hFF;
            15'd7553: data <= 8'hFF;
            15'd7554: data <= 8'hFF;
            15'd7555: data <= 8'h80;
            15'd7556: data <= 8'h00;
            15'd7557: data <= 8'h00;
            15'd7558: data <= 8'h00;
            15'd7559: data <= 8'h00;
            15'd7560: data <= 8'h00;
            15'd7561: data <= 8'h00;
            15'd7562: data <= 8'h00;
            15'd7563: data <= 8'h00;
            15'd7564: data <= 8'h01;
            15'd7565: data <= 8'hFF;
            15'd7566: data <= 8'hFF;
            15'd7567: data <= 8'hFF;
            15'd7568: data <= 8'hFF;
            15'd7569: data <= 8'hFF;
            15'd7570: data <= 8'hFF;
            15'd7571: data <= 8'h9C;
            15'd7572: data <= 8'h3F;
            15'd7573: data <= 8'hFF;
            15'd7574: data <= 8'hFF;
            15'd7575: data <= 8'hFF;
            15'd7576: data <= 8'hFF;
            15'd7577: data <= 8'hFF;
            15'd7578: data <= 8'hF0;
            15'd7579: data <= 8'hF1;
            15'd7580: data <= 8'hFF;
            15'd7581: data <= 8'hFF;
            15'd7582: data <= 8'hFF;
            15'd7583: data <= 8'hFF;
            15'd7584: data <= 8'hFF;
            15'd7585: data <= 8'h80;
            15'd7586: data <= 8'h00;
            15'd7587: data <= 8'h00;
            15'd7588: data <= 8'h00;
            15'd7589: data <= 8'h00;
            15'd7590: data <= 8'h00;
            15'd7591: data <= 8'h00;
            15'd7592: data <= 8'h00;
            15'd7593: data <= 8'h00;
            15'd7594: data <= 8'h01;
            15'd7595: data <= 8'hFF;
            15'd7596: data <= 8'hFF;
            15'd7597: data <= 8'hFF;
            15'd7598: data <= 8'hFF;
            15'd7599: data <= 8'hFF;
            15'd7600: data <= 8'hFF;
            15'd7601: data <= 8'h0C;
            15'd7602: data <= 8'h1F;
            15'd7603: data <= 8'hFF;
            15'd7604: data <= 8'hFE;
            15'd7605: data <= 8'h07;
            15'd7606: data <= 8'hFF;
            15'd7607: data <= 8'hFF;
            15'd7608: data <= 8'hE1;
            15'd7609: data <= 8'hE1;
            15'd7610: data <= 8'hFF;
            15'd7611: data <= 8'hFF;
            15'd7612: data <= 8'hFF;
            15'd7613: data <= 8'hFF;
            15'd7614: data <= 8'hFF;
            15'd7615: data <= 8'h80;
            15'd7616: data <= 8'h00;
            15'd7617: data <= 8'h00;
            15'd7618: data <= 8'h00;
            15'd7619: data <= 8'h00;
            15'd7620: data <= 8'h00;
            15'd7621: data <= 8'h00;
            15'd7622: data <= 8'h00;
            15'd7623: data <= 8'h00;
            15'd7624: data <= 8'h01;
            15'd7625: data <= 8'hFF;
            15'd7626: data <= 8'hFF;
            15'd7627: data <= 8'hFF;
            15'd7628: data <= 8'hFF;
            15'd7629: data <= 8'hFF;
            15'd7630: data <= 8'hFE;
            15'd7631: data <= 8'h0C;
            15'd7632: data <= 8'h3F;
            15'd7633: data <= 8'hFF;
            15'd7634: data <= 8'hF8;
            15'd7635: data <= 8'h01;
            15'd7636: data <= 8'hFF;
            15'd7637: data <= 8'hFF;
            15'd7638: data <= 8'hE1;
            15'd7639: data <= 8'hE1;
            15'd7640: data <= 8'hFF;
            15'd7641: data <= 8'hFF;
            15'd7642: data <= 8'hFF;
            15'd7643: data <= 8'hFF;
            15'd7644: data <= 8'hFF;
            15'd7645: data <= 8'h80;
            15'd7646: data <= 8'h00;
            15'd7647: data <= 8'h00;
            15'd7648: data <= 8'h00;
            15'd7649: data <= 8'h00;
            15'd7650: data <= 8'h00;
            15'd7651: data <= 8'h00;
            15'd7652: data <= 8'h00;
            15'd7653: data <= 8'h00;
            15'd7654: data <= 8'h01;
            15'd7655: data <= 8'hFF;
            15'd7656: data <= 8'hFF;
            15'd7657: data <= 8'hFF;
            15'd7658: data <= 8'hFF;
            15'd7659: data <= 8'hFF;
            15'd7660: data <= 8'hFE;
            15'd7661: data <= 8'h1C;
            15'd7662: data <= 8'h3F;
            15'd7663: data <= 8'hFF;
            15'd7664: data <= 8'hF0;
            15'd7665: data <= 8'h00;
            15'd7666: data <= 8'hFF;
            15'd7667: data <= 8'hFF;
            15'd7668: data <= 8'hF1;
            15'd7669: data <= 8'hF1;
            15'd7670: data <= 8'hFF;
            15'd7671: data <= 8'hFF;
            15'd7672: data <= 8'hFF;
            15'd7673: data <= 8'hFF;
            15'd7674: data <= 8'hFF;
            15'd7675: data <= 8'h80;
            15'd7676: data <= 8'h00;
            15'd7677: data <= 8'h00;
            15'd7678: data <= 8'h00;
            15'd7679: data <= 8'h00;
            15'd7680: data <= 8'h00;
            15'd7681: data <= 8'h00;
            15'd7682: data <= 8'h00;
            15'd7683: data <= 8'h00;
            15'd7684: data <= 8'h01;
            15'd7685: data <= 8'hFF;
            15'd7686: data <= 8'hFF;
            15'd7687: data <= 8'hFF;
            15'd7688: data <= 8'hFF;
            15'd7689: data <= 8'hFF;
            15'd7690: data <= 8'hFE;
            15'd7691: data <= 8'h1C;
            15'd7692: data <= 8'h7F;
            15'd7693: data <= 8'hFF;
            15'd7694: data <= 8'hE0;
            15'd7695: data <= 8'h00;
            15'd7696: data <= 8'h7F;
            15'd7697: data <= 8'hFF;
            15'd7698: data <= 8'hF3;
            15'd7699: data <= 8'hF3;
            15'd7700: data <= 8'hFF;
            15'd7701: data <= 8'hFF;
            15'd7702: data <= 8'hFF;
            15'd7703: data <= 8'hFF;
            15'd7704: data <= 8'hFF;
            15'd7705: data <= 8'h80;
            15'd7706: data <= 8'h00;
            15'd7707: data <= 8'h00;
            15'd7708: data <= 8'h00;
            15'd7709: data <= 8'h00;
            15'd7710: data <= 8'h00;
            15'd7711: data <= 8'h00;
            15'd7712: data <= 8'h00;
            15'd7713: data <= 8'h00;
            15'd7714: data <= 8'h01;
            15'd7715: data <= 8'hFF;
            15'd7716: data <= 8'hFF;
            15'd7717: data <= 8'hFF;
            15'd7718: data <= 8'hFF;
            15'd7719: data <= 8'hFF;
            15'd7720: data <= 8'hFF;
            15'd7721: data <= 8'h1C;
            15'd7722: data <= 8'hFF;
            15'd7723: data <= 8'hFF;
            15'd7724: data <= 8'hC0;
            15'd7725: data <= 8'h40;
            15'd7726: data <= 8'h3F;
            15'd7727: data <= 8'hF8;
            15'd7728: data <= 8'hFF;
            15'd7729: data <= 8'hFF;
            15'd7730: data <= 8'hFF;
            15'd7731: data <= 8'hFF;
            15'd7732: data <= 8'hFF;
            15'd7733: data <= 8'hFF;
            15'd7734: data <= 8'hFF;
            15'd7735: data <= 8'h80;
            15'd7736: data <= 8'h00;
            15'd7737: data <= 8'h00;
            15'd7738: data <= 8'h00;
            15'd7739: data <= 8'h00;
            15'd7740: data <= 8'h00;
            15'd7741: data <= 8'h00;
            15'd7742: data <= 8'h00;
            15'd7743: data <= 8'h00;
            15'd7744: data <= 8'h01;
            15'd7745: data <= 8'hFF;
            15'd7746: data <= 8'hFF;
            15'd7747: data <= 8'hFF;
            15'd7748: data <= 8'hFF;
            15'd7749: data <= 8'hFF;
            15'd7750: data <= 8'hFF;
            15'd7751: data <= 8'hBF;
            15'd7752: data <= 8'hFF;
            15'd7753: data <= 8'hFF;
            15'd7754: data <= 8'h81;
            15'd7755: data <= 8'hF0;
            15'd7756: data <= 8'h1F;
            15'd7757: data <= 8'hF8;
            15'd7758: data <= 8'h7F;
            15'd7759: data <= 8'hFF;
            15'd7760: data <= 8'hFF;
            15'd7761: data <= 8'hFF;
            15'd7762: data <= 8'hFF;
            15'd7763: data <= 8'hFF;
            15'd7764: data <= 8'hFF;
            15'd7765: data <= 8'h80;
            15'd7766: data <= 8'h00;
            15'd7767: data <= 8'h00;
            15'd7768: data <= 8'h00;
            15'd7769: data <= 8'h00;
            15'd7770: data <= 8'h00;
            15'd7771: data <= 8'h00;
            15'd7772: data <= 8'h00;
            15'd7773: data <= 8'h00;
            15'd7774: data <= 8'h01;
            15'd7775: data <= 8'hFF;
            15'd7776: data <= 8'hFF;
            15'd7777: data <= 8'hFF;
            15'd7778: data <= 8'hFF;
            15'd7779: data <= 8'hFF;
            15'd7780: data <= 8'hFF;
            15'd7781: data <= 8'hFF;
            15'd7782: data <= 8'hFF;
            15'd7783: data <= 8'hFF;
            15'd7784: data <= 8'h83;
            15'd7785: data <= 8'hFC;
            15'd7786: data <= 8'h1F;
            15'd7787: data <= 8'hF0;
            15'd7788: data <= 8'h7F;
            15'd7789: data <= 8'hFF;
            15'd7790: data <= 8'hFF;
            15'd7791: data <= 8'hFF;
            15'd7792: data <= 8'hFF;
            15'd7793: data <= 8'hFF;
            15'd7794: data <= 8'hFF;
            15'd7795: data <= 8'h80;
            15'd7796: data <= 8'h00;
            15'd7797: data <= 8'h00;
            15'd7798: data <= 8'h00;
            15'd7799: data <= 8'h00;
            15'd7800: data <= 8'h00;
            15'd7801: data <= 8'h00;
            15'd7802: data <= 8'h00;
            15'd7803: data <= 8'h00;
            15'd7804: data <= 8'h01;
            15'd7805: data <= 8'hFF;
            15'd7806: data <= 8'hFF;
            15'd7807: data <= 8'hFF;
            15'd7808: data <= 8'hFF;
            15'd7809: data <= 8'hFF;
            15'd7810: data <= 8'hFF;
            15'd7811: data <= 8'hFF;
            15'd7812: data <= 8'hFF;
            15'd7813: data <= 8'hFF;
            15'd7814: data <= 8'h07;
            15'd7815: data <= 8'hFE;
            15'd7816: data <= 8'h1F;
            15'd7817: data <= 8'hE0;
            15'd7818: data <= 8'hFF;
            15'd7819: data <= 8'hFF;
            15'd7820: data <= 8'hFF;
            15'd7821: data <= 8'hFF;
            15'd7822: data <= 8'hFF;
            15'd7823: data <= 8'hFF;
            15'd7824: data <= 8'hFF;
            15'd7825: data <= 8'h80;
            15'd7826: data <= 8'h00;
            15'd7827: data <= 8'h00;
            15'd7828: data <= 8'h00;
            15'd7829: data <= 8'h00;
            15'd7830: data <= 8'h00;
            15'd7831: data <= 8'h00;
            15'd7832: data <= 8'h00;
            15'd7833: data <= 8'h00;
            15'd7834: data <= 8'h01;
            15'd7835: data <= 8'hFF;
            15'd7836: data <= 8'hFF;
            15'd7837: data <= 8'hFF;
            15'd7838: data <= 8'hFF;
            15'd7839: data <= 8'hFF;
            15'd7840: data <= 8'hFF;
            15'd7841: data <= 8'hFF;
            15'd7842: data <= 8'hFF;
            15'd7843: data <= 8'hFF;
            15'd7844: data <= 8'h0F;
            15'd7845: data <= 8'hFF;
            15'd7846: data <= 8'hFF;
            15'd7847: data <= 8'hE0;
            15'd7848: data <= 8'hFF;
            15'd7849: data <= 8'hFF;
            15'd7850: data <= 8'hFF;
            15'd7851: data <= 8'hFF;
            15'd7852: data <= 8'hFF;
            15'd7853: data <= 8'hFF;
            15'd7854: data <= 8'hFF;
            15'd7855: data <= 8'h80;
            15'd7856: data <= 8'h00;
            15'd7857: data <= 8'h00;
            15'd7858: data <= 8'h00;
            15'd7859: data <= 8'h00;
            15'd7860: data <= 8'h00;
            15'd7861: data <= 8'h00;
            15'd7862: data <= 8'h00;
            15'd7863: data <= 8'h00;
            15'd7864: data <= 8'h01;
            15'd7865: data <= 8'hFF;
            15'd7866: data <= 8'hFF;
            15'd7867: data <= 8'hFF;
            15'd7868: data <= 8'hFF;
            15'd7869: data <= 8'hFF;
            15'd7870: data <= 8'hFF;
            15'd7871: data <= 8'hFF;
            15'd7872: data <= 8'hFF;
            15'd7873: data <= 8'hFF;
            15'd7874: data <= 8'h9F;
            15'd7875: data <= 8'hFF;
            15'd7876: data <= 8'hFF;
            15'd7877: data <= 8'hC1;
            15'd7878: data <= 8'hFF;
            15'd7879: data <= 8'hFF;
            15'd7880: data <= 8'hFF;
            15'd7881: data <= 8'hFF;
            15'd7882: data <= 8'hFF;
            15'd7883: data <= 8'hFF;
            15'd7884: data <= 8'hFF;
            15'd7885: data <= 8'h80;
            15'd7886: data <= 8'h00;
            15'd7887: data <= 8'h00;
            15'd7888: data <= 8'h00;
            15'd7889: data <= 8'h00;
            15'd7890: data <= 8'h00;
            15'd7891: data <= 8'h00;
            15'd7892: data <= 8'h00;
            15'd7893: data <= 8'h00;
            15'd7894: data <= 8'h01;
            15'd7895: data <= 8'hFF;
            15'd7896: data <= 8'hFF;
            15'd7897: data <= 8'hFF;
            15'd7898: data <= 8'hFF;
            15'd7899: data <= 8'hFF;
            15'd7900: data <= 8'hFF;
            15'd7901: data <= 8'hFF;
            15'd7902: data <= 8'hFF;
            15'd7903: data <= 8'hFF;
            15'd7904: data <= 8'hFF;
            15'd7905: data <= 8'hFF;
            15'd7906: data <= 8'hFF;
            15'd7907: data <= 8'hC3;
            15'd7908: data <= 8'hFF;
            15'd7909: data <= 8'hFF;
            15'd7910: data <= 8'hFF;
            15'd7911: data <= 8'hFF;
            15'd7912: data <= 8'hFF;
            15'd7913: data <= 8'hFF;
            15'd7914: data <= 8'hFF;
            15'd7915: data <= 8'h80;
            15'd7916: data <= 8'h00;
            15'd7917: data <= 8'h00;
            15'd7918: data <= 8'h00;
            15'd7919: data <= 8'h00;
            15'd7920: data <= 8'h00;
            15'd7921: data <= 8'h00;
            15'd7922: data <= 8'h00;
            15'd7923: data <= 8'h00;
            15'd7924: data <= 8'h01;
            15'd7925: data <= 8'hFF;
            15'd7926: data <= 8'hFF;
            15'd7927: data <= 8'hFF;
            15'd7928: data <= 8'hFF;
            15'd7929: data <= 8'hFF;
            15'd7930: data <= 8'hFF;
            15'd7931: data <= 8'hFF;
            15'd7932: data <= 8'hFF;
            15'd7933: data <= 8'hFF;
            15'd7934: data <= 8'hFF;
            15'd7935: data <= 8'hFF;
            15'd7936: data <= 8'hFF;
            15'd7937: data <= 8'h83;
            15'd7938: data <= 8'hFF;
            15'd7939: data <= 8'hFF;
            15'd7940: data <= 8'hFF;
            15'd7941: data <= 8'hFF;
            15'd7942: data <= 8'hFF;
            15'd7943: data <= 8'hFF;
            15'd7944: data <= 8'hFF;
            15'd7945: data <= 8'h80;
            15'd7946: data <= 8'h00;
            15'd7947: data <= 8'h00;
            15'd7948: data <= 8'h00;
            15'd7949: data <= 8'h00;
            15'd7950: data <= 8'h00;
            15'd7951: data <= 8'h00;
            15'd7952: data <= 8'h00;
            15'd7953: data <= 8'h00;
            15'd7954: data <= 8'h01;
            15'd7955: data <= 8'hFF;
            15'd7956: data <= 8'hFF;
            15'd7957: data <= 8'hFF;
            15'd7958: data <= 8'hFF;
            15'd7959: data <= 8'hFF;
            15'd7960: data <= 8'hFF;
            15'd7961: data <= 8'hFF;
            15'd7962: data <= 8'hFF;
            15'd7963: data <= 8'hFF;
            15'd7964: data <= 8'hFF;
            15'd7965: data <= 8'hFF;
            15'd7966: data <= 8'hFF;
            15'd7967: data <= 8'h87;
            15'd7968: data <= 8'hFF;
            15'd7969: data <= 8'h1F;
            15'd7970: data <= 8'hFF;
            15'd7971: data <= 8'hFF;
            15'd7972: data <= 8'hFF;
            15'd7973: data <= 8'hFF;
            15'd7974: data <= 8'hFF;
            15'd7975: data <= 8'h80;
            15'd7976: data <= 8'h00;
            15'd7977: data <= 8'h00;
            15'd7978: data <= 8'h00;
            15'd7979: data <= 8'h00;
            15'd7980: data <= 8'h00;
            15'd7981: data <= 8'h00;
            15'd7982: data <= 8'h00;
            15'd7983: data <= 8'h00;
            15'd7984: data <= 8'h01;
            15'd7985: data <= 8'hFF;
            15'd7986: data <= 8'hFF;
            15'd7987: data <= 8'hFF;
            15'd7988: data <= 8'hFF;
            15'd7989: data <= 8'hFF;
            15'd7990: data <= 8'hFF;
            15'd7991: data <= 8'hFF;
            15'd7992: data <= 8'hFF;
            15'd7993: data <= 8'hFF;
            15'd7994: data <= 8'hFF;
            15'd7995: data <= 8'hFF;
            15'd7996: data <= 8'hFF;
            15'd7997: data <= 8'h07;
            15'd7998: data <= 8'hFE;
            15'd7999: data <= 8'h1F;
            15'd8000: data <= 8'hFF;
            15'd8001: data <= 8'hFF;
            15'd8002: data <= 8'hFF;
            15'd8003: data <= 8'hFF;
            15'd8004: data <= 8'hFF;
            15'd8005: data <= 8'h80;
            15'd8006: data <= 8'h00;
            15'd8007: data <= 8'h00;
            15'd8008: data <= 8'h00;
            15'd8009: data <= 8'h00;
            15'd8010: data <= 8'h00;
            15'd8011: data <= 8'h00;
            15'd8012: data <= 8'h00;
            15'd8013: data <= 8'h00;
            15'd8014: data <= 8'h01;
            15'd8015: data <= 8'hFF;
            15'd8016: data <= 8'hFF;
            15'd8017: data <= 8'hFF;
            15'd8018: data <= 8'hFF;
            15'd8019: data <= 8'hFF;
            15'd8020: data <= 8'hFF;
            15'd8021: data <= 8'hFF;
            15'd8022: data <= 8'hFF;
            15'd8023: data <= 8'hFF;
            15'd8024: data <= 8'hFF;
            15'd8025: data <= 8'hFF;
            15'd8026: data <= 8'hFE;
            15'd8027: data <= 8'h0F;
            15'd8028: data <= 8'hFC;
            15'd8029: data <= 8'h1F;
            15'd8030: data <= 8'hFF;
            15'd8031: data <= 8'hFF;
            15'd8032: data <= 8'hFF;
            15'd8033: data <= 8'hFF;
            15'd8034: data <= 8'hFF;
            15'd8035: data <= 8'h80;
            15'd8036: data <= 8'h00;
            15'd8037: data <= 8'h00;
            15'd8038: data <= 8'h00;
            15'd8039: data <= 8'h00;
            15'd8040: data <= 8'h00;
            15'd8041: data <= 8'h00;
            15'd8042: data <= 8'h00;
            15'd8043: data <= 8'h00;
            15'd8044: data <= 8'h01;
            15'd8045: data <= 8'hFF;
            15'd8046: data <= 8'hFF;
            15'd8047: data <= 8'hFF;
            15'd8048: data <= 8'hFF;
            15'd8049: data <= 8'hFF;
            15'd8050: data <= 8'hFF;
            15'd8051: data <= 8'hFF;
            15'd8052: data <= 8'hFF;
            15'd8053: data <= 8'hFF;
            15'd8054: data <= 8'hFF;
            15'd8055: data <= 8'hFF;
            15'd8056: data <= 8'hFE;
            15'd8057: data <= 8'h0F;
            15'd8058: data <= 8'hF8;
            15'd8059: data <= 8'h3F;
            15'd8060: data <= 8'hFF;
            15'd8061: data <= 8'hFF;
            15'd8062: data <= 8'hFF;
            15'd8063: data <= 8'hFF;
            15'd8064: data <= 8'hFF;
            15'd8065: data <= 8'h80;
            15'd8066: data <= 8'h00;
            15'd8067: data <= 8'h00;
            15'd8068: data <= 8'h00;
            15'd8069: data <= 8'h00;
            15'd8070: data <= 8'h00;
            15'd8071: data <= 8'h00;
            15'd8072: data <= 8'h00;
            15'd8073: data <= 8'h00;
            15'd8074: data <= 8'h01;
            15'd8075: data <= 8'hFF;
            15'd8076: data <= 8'hFF;
            15'd8077: data <= 8'hFF;
            15'd8078: data <= 8'hFF;
            15'd8079: data <= 8'hFF;
            15'd8080: data <= 8'hFF;
            15'd8081: data <= 8'hFF;
            15'd8082: data <= 8'hFF;
            15'd8083: data <= 8'hFF;
            15'd8084: data <= 8'hFF;
            15'd8085: data <= 8'hFF;
            15'd8086: data <= 8'hFE;
            15'd8087: data <= 8'h1F;
            15'd8088: data <= 8'hF8;
            15'd8089: data <= 8'h3F;
            15'd8090: data <= 8'hFF;
            15'd8091: data <= 8'hFF;
            15'd8092: data <= 8'hFF;
            15'd8093: data <= 8'hFF;
            15'd8094: data <= 8'hFF;
            15'd8095: data <= 8'h80;
            15'd8096: data <= 8'h00;
            15'd8097: data <= 8'h00;
            15'd8098: data <= 8'h00;
            15'd8099: data <= 8'h00;
            15'd8100: data <= 8'h00;
            15'd8101: data <= 8'h00;
            15'd8102: data <= 8'h00;
            15'd8103: data <= 8'h00;
            15'd8104: data <= 8'h01;
            15'd8105: data <= 8'hFF;
            15'd8106: data <= 8'hFF;
            15'd8107: data <= 8'hFF;
            15'd8108: data <= 8'hFF;
            15'd8109: data <= 8'hFF;
            15'd8110: data <= 8'hFF;
            15'd8111: data <= 8'hFF;
            15'd8112: data <= 8'hFF;
            15'd8113: data <= 8'hFF;
            15'd8114: data <= 8'hFF;
            15'd8115: data <= 8'hFF;
            15'd8116: data <= 8'hFC;
            15'd8117: data <= 8'h1F;
            15'd8118: data <= 8'hF0;
            15'd8119: data <= 8'h7F;
            15'd8120: data <= 8'hFF;
            15'd8121: data <= 8'hFF;
            15'd8122: data <= 8'hFF;
            15'd8123: data <= 8'hFF;
            15'd8124: data <= 8'hFF;
            15'd8125: data <= 8'h80;
            15'd8126: data <= 8'h00;
            15'd8127: data <= 8'h00;
            15'd8128: data <= 8'h00;
            15'd8129: data <= 8'h00;
            15'd8130: data <= 8'h00;
            15'd8131: data <= 8'h00;
            15'd8132: data <= 8'h00;
            15'd8133: data <= 8'h00;
            15'd8134: data <= 8'h01;
            15'd8135: data <= 8'hFF;
            15'd8136: data <= 8'hFF;
            15'd8137: data <= 8'hFF;
            15'd8138: data <= 8'hFF;
            15'd8139: data <= 8'hFF;
            15'd8140: data <= 8'hFF;
            15'd8141: data <= 8'hFF;
            15'd8142: data <= 8'hFF;
            15'd8143: data <= 8'hFF;
            15'd8144: data <= 8'hFF;
            15'd8145: data <= 8'hFF;
            15'd8146: data <= 8'hFC;
            15'd8147: data <= 8'h3F;
            15'd8148: data <= 8'hE0;
            15'd8149: data <= 8'hFF;
            15'd8150: data <= 8'hFF;
            15'd8151: data <= 8'hFF;
            15'd8152: data <= 8'hFF;
            15'd8153: data <= 8'hFF;
            15'd8154: data <= 8'hFF;
            15'd8155: data <= 8'h80;
            15'd8156: data <= 8'h00;
            15'd8157: data <= 8'h00;
            15'd8158: data <= 8'h00;
            15'd8159: data <= 8'h00;
            15'd8160: data <= 8'h00;
            15'd8161: data <= 8'h00;
            15'd8162: data <= 8'h00;
            15'd8163: data <= 8'h00;
            15'd8164: data <= 8'h01;
            15'd8165: data <= 8'hFF;
            15'd8166: data <= 8'hFF;
            15'd8167: data <= 8'hFF;
            15'd8168: data <= 8'hFF;
            15'd8169: data <= 8'hFF;
            15'd8170: data <= 8'hFF;
            15'd8171: data <= 8'hFF;
            15'd8172: data <= 8'hFF;
            15'd8173: data <= 8'hFF;
            15'd8174: data <= 8'hFF;
            15'd8175: data <= 8'hFF;
            15'd8176: data <= 8'hFC;
            15'd8177: data <= 8'h3F;
            15'd8178: data <= 8'hC0;
            15'd8179: data <= 8'hFF;
            15'd8180: data <= 8'hFF;
            15'd8181: data <= 8'hFF;
            15'd8182: data <= 8'hFF;
            15'd8183: data <= 8'hFF;
            15'd8184: data <= 8'hFF;
            15'd8185: data <= 8'h80;
            15'd8186: data <= 8'h00;
            15'd8187: data <= 8'h00;
            15'd8188: data <= 8'h00;
            15'd8189: data <= 8'h00;
            15'd8190: data <= 8'h00;
            15'd8191: data <= 8'h00;
            15'd8192: data <= 8'h00;
            15'd8193: data <= 8'h00;
            15'd8194: data <= 8'h01;
            15'd8195: data <= 8'hFF;
            15'd8196: data <= 8'hFF;
            15'd8197: data <= 8'hFF;
            15'd8198: data <= 8'hFF;
            15'd8199: data <= 8'hFF;
            15'd8200: data <= 8'hFF;
            15'd8201: data <= 8'hFF;
            15'd8202: data <= 8'hFF;
            15'd8203: data <= 8'hFF;
            15'd8204: data <= 8'hFF;
            15'd8205: data <= 8'hFF;
            15'd8206: data <= 8'hF8;
            15'd8207: data <= 8'h7F;
            15'd8208: data <= 8'h81;
            15'd8209: data <= 8'hFF;
            15'd8210: data <= 8'hFF;
            15'd8211: data <= 8'hFF;
            15'd8212: data <= 8'hFF;
            15'd8213: data <= 8'hFF;
            15'd8214: data <= 8'hFF;
            15'd8215: data <= 8'h80;
            15'd8216: data <= 8'h00;
            15'd8217: data <= 8'h00;
            15'd8218: data <= 8'h00;
            15'd8219: data <= 8'h00;
            15'd8220: data <= 8'h00;
            15'd8221: data <= 8'h00;
            15'd8222: data <= 8'h00;
            15'd8223: data <= 8'h00;
            15'd8224: data <= 8'h01;
            15'd8225: data <= 8'hFF;
            15'd8226: data <= 8'hFF;
            15'd8227: data <= 8'hFF;
            15'd8228: data <= 8'hFF;
            15'd8229: data <= 8'hFF;
            15'd8230: data <= 8'hFF;
            15'd8231: data <= 8'hFF;
            15'd8232: data <= 8'hFF;
            15'd8233: data <= 8'hFF;
            15'd8234: data <= 8'hFF;
            15'd8235: data <= 8'hFF;
            15'd8236: data <= 8'hF8;
            15'd8237: data <= 8'h7F;
            15'd8238: data <= 8'h03;
            15'd8239: data <= 8'hFF;
            15'd8240: data <= 8'hFF;
            15'd8241: data <= 8'hFF;
            15'd8242: data <= 8'hFF;
            15'd8243: data <= 8'hFF;
            15'd8244: data <= 8'hFF;
            15'd8245: data <= 8'h80;
            15'd8246: data <= 8'h00;
            15'd8247: data <= 8'h00;
            15'd8248: data <= 8'h00;
            15'd8249: data <= 8'h00;
            15'd8250: data <= 8'h00;
            15'd8251: data <= 8'h00;
            15'd8252: data <= 8'h00;
            15'd8253: data <= 8'h00;
            15'd8254: data <= 8'h01;
            15'd8255: data <= 8'hFF;
            15'd8256: data <= 8'hFF;
            15'd8257: data <= 8'hFF;
            15'd8258: data <= 8'hFF;
            15'd8259: data <= 8'hFF;
            15'd8260: data <= 8'hFF;
            15'd8261: data <= 8'hFF;
            15'd8262: data <= 8'hFF;
            15'd8263: data <= 8'hFF;
            15'd8264: data <= 8'hFF;
            15'd8265: data <= 8'hFF;
            15'd8266: data <= 8'hF8;
            15'd8267: data <= 8'h7E;
            15'd8268: data <= 8'h07;
            15'd8269: data <= 8'hFF;
            15'd8270: data <= 8'hFF;
            15'd8271: data <= 8'hFF;
            15'd8272: data <= 8'hFF;
            15'd8273: data <= 8'hFF;
            15'd8274: data <= 8'hFF;
            15'd8275: data <= 8'h80;
            15'd8276: data <= 8'h00;
            15'd8277: data <= 8'h00;
            15'd8278: data <= 8'h00;
            15'd8279: data <= 8'h00;
            15'd8280: data <= 8'h00;
            15'd8281: data <= 8'h00;
            15'd8282: data <= 8'h00;
            15'd8283: data <= 8'h00;
            15'd8284: data <= 8'h01;
            15'd8285: data <= 8'hFF;
            15'd8286: data <= 8'hFF;
            15'd8287: data <= 8'hFF;
            15'd8288: data <= 8'hFF;
            15'd8289: data <= 8'hFF;
            15'd8290: data <= 8'hFF;
            15'd8291: data <= 8'hFF;
            15'd8292: data <= 8'hFF;
            15'd8293: data <= 8'hFF;
            15'd8294: data <= 8'hFF;
            15'd8295: data <= 8'hFF;
            15'd8296: data <= 8'hF8;
            15'd8297: data <= 8'h7C;
            15'd8298: data <= 8'h0F;
            15'd8299: data <= 8'hFF;
            15'd8300: data <= 8'hFF;
            15'd8301: data <= 8'hFF;
            15'd8302: data <= 8'hFF;
            15'd8303: data <= 8'hFF;
            15'd8304: data <= 8'hFF;
            15'd8305: data <= 8'h80;
            15'd8306: data <= 8'h00;
            15'd8307: data <= 8'h00;
            15'd8308: data <= 8'h00;
            15'd8309: data <= 8'h00;
            15'd8310: data <= 8'h00;
            15'd8311: data <= 8'h00;
            15'd8312: data <= 8'h00;
            15'd8313: data <= 8'h00;
            15'd8314: data <= 8'h01;
            15'd8315: data <= 8'hFF;
            15'd8316: data <= 8'hFF;
            15'd8317: data <= 8'hFF;
            15'd8318: data <= 8'hFF;
            15'd8319: data <= 8'hFF;
            15'd8320: data <= 8'hFF;
            15'd8321: data <= 8'hFF;
            15'd8322: data <= 8'hFF;
            15'd8323: data <= 8'hFF;
            15'd8324: data <= 8'hFF;
            15'd8325: data <= 8'hFF;
            15'd8326: data <= 8'hF8;
            15'd8327: data <= 8'h70;
            15'd8328: data <= 8'h1F;
            15'd8329: data <= 8'hFF;
            15'd8330: data <= 8'hFF;
            15'd8331: data <= 8'hFF;
            15'd8332: data <= 8'hFF;
            15'd8333: data <= 8'hFF;
            15'd8334: data <= 8'hFF;
            15'd8335: data <= 8'h80;
            15'd8336: data <= 8'h00;
            15'd8337: data <= 8'h00;
            15'd8338: data <= 8'h00;
            15'd8339: data <= 8'h00;
            15'd8340: data <= 8'h00;
            15'd8341: data <= 8'h00;
            15'd8342: data <= 8'h00;
            15'd8343: data <= 8'h00;
            15'd8344: data <= 8'h01;
            15'd8345: data <= 8'hFF;
            15'd8346: data <= 8'hFF;
            15'd8347: data <= 8'hFF;
            15'd8348: data <= 8'hFF;
            15'd8349: data <= 8'hFF;
            15'd8350: data <= 8'hFF;
            15'd8351: data <= 8'hFF;
            15'd8352: data <= 8'hFF;
            15'd8353: data <= 8'hFF;
            15'd8354: data <= 8'hFF;
            15'd8355: data <= 8'hFF;
            15'd8356: data <= 8'hF8;
            15'd8357: data <= 8'h40;
            15'd8358: data <= 8'h3F;
            15'd8359: data <= 8'hFF;
            15'd8360: data <= 8'hFF;
            15'd8361: data <= 8'hFF;
            15'd8362: data <= 8'hFF;
            15'd8363: data <= 8'hFF;
            15'd8364: data <= 8'hFF;
            15'd8365: data <= 8'h80;
            15'd8366: data <= 8'h00;
            15'd8367: data <= 8'h00;
            15'd8368: data <= 8'h00;
            15'd8369: data <= 8'h00;
            15'd8370: data <= 8'h00;
            15'd8371: data <= 8'h00;
            15'd8372: data <= 8'h00;
            15'd8373: data <= 8'h00;
            15'd8374: data <= 8'h01;
            15'd8375: data <= 8'hFF;
            15'd8376: data <= 8'hFF;
            15'd8377: data <= 8'hFF;
            15'd8378: data <= 8'hFF;
            15'd8379: data <= 8'hFF;
            15'd8380: data <= 8'hFF;
            15'd8381: data <= 8'hFF;
            15'd8382: data <= 8'hFF;
            15'd8383: data <= 8'hFF;
            15'd8384: data <= 8'hFF;
            15'd8385: data <= 8'hFF;
            15'd8386: data <= 8'hF8;
            15'd8387: data <= 8'h00;
            15'd8388: data <= 8'h7F;
            15'd8389: data <= 8'hFF;
            15'd8390: data <= 8'hFF;
            15'd8391: data <= 8'hFF;
            15'd8392: data <= 8'hFF;
            15'd8393: data <= 8'hFF;
            15'd8394: data <= 8'hFF;
            15'd8395: data <= 8'h80;
            15'd8396: data <= 8'h00;
            15'd8397: data <= 8'h00;
            15'd8398: data <= 8'h00;
            15'd8399: data <= 8'h00;
            15'd8400: data <= 8'h00;
            15'd8401: data <= 8'h00;
            15'd8402: data <= 8'h00;
            15'd8403: data <= 8'h00;
            15'd8404: data <= 8'h01;
            15'd8405: data <= 8'hFF;
            15'd8406: data <= 8'hFF;
            15'd8407: data <= 8'hFF;
            15'd8408: data <= 8'hFF;
            15'd8409: data <= 8'hFF;
            15'd8410: data <= 8'hFF;
            15'd8411: data <= 8'hFF;
            15'd8412: data <= 8'hFF;
            15'd8413: data <= 8'hFF;
            15'd8414: data <= 8'hFF;
            15'd8415: data <= 8'hFF;
            15'd8416: data <= 8'hFC;
            15'd8417: data <= 8'h00;
            15'd8418: data <= 8'hFF;
            15'd8419: data <= 8'hFF;
            15'd8420: data <= 8'hFF;
            15'd8421: data <= 8'hFF;
            15'd8422: data <= 8'hFF;
            15'd8423: data <= 8'hFF;
            15'd8424: data <= 8'hFF;
            15'd8425: data <= 8'h80;
            15'd8426: data <= 8'h00;
            15'd8427: data <= 8'h00;
            15'd8428: data <= 8'h00;
            15'd8429: data <= 8'h00;
            15'd8430: data <= 8'h00;
            15'd8431: data <= 8'h00;
            15'd8432: data <= 8'h00;
            15'd8433: data <= 8'h00;
            15'd8434: data <= 8'h01;
            15'd8435: data <= 8'hFF;
            15'd8436: data <= 8'hFF;
            15'd8437: data <= 8'hFF;
            15'd8438: data <= 8'hFF;
            15'd8439: data <= 8'hFF;
            15'd8440: data <= 8'hFF;
            15'd8441: data <= 8'hFF;
            15'd8442: data <= 8'hFF;
            15'd8443: data <= 8'hFF;
            15'd8444: data <= 8'hFF;
            15'd8445: data <= 8'hCF;
            15'd8446: data <= 8'hFC;
            15'd8447: data <= 8'h03;
            15'd8448: data <= 8'hFF;
            15'd8449: data <= 8'hFF;
            15'd8450: data <= 8'hFF;
            15'd8451: data <= 8'hFF;
            15'd8452: data <= 8'hFF;
            15'd8453: data <= 8'hFF;
            15'd8454: data <= 8'hFF;
            15'd8455: data <= 8'h80;
            15'd8456: data <= 8'h00;
            15'd8457: data <= 8'h00;
            15'd8458: data <= 8'h00;
            15'd8459: data <= 8'h00;
            15'd8460: data <= 8'h00;
            15'd8461: data <= 8'h00;
            15'd8462: data <= 8'h00;
            15'd8463: data <= 8'h00;
            15'd8464: data <= 8'h01;
            15'd8465: data <= 8'hFF;
            15'd8466: data <= 8'hFF;
            15'd8467: data <= 8'hFF;
            15'd8468: data <= 8'hFF;
            15'd8469: data <= 8'hFF;
            15'd8470: data <= 8'hFF;
            15'd8471: data <= 8'hFF;
            15'd8472: data <= 8'hFF;
            15'd8473: data <= 8'hFF;
            15'd8474: data <= 8'hFF;
            15'd8475: data <= 8'h8F;
            15'd8476: data <= 8'hFF;
            15'd8477: data <= 8'h0F;
            15'd8478: data <= 8'hFF;
            15'd8479: data <= 8'hFF;
            15'd8480: data <= 8'hFF;
            15'd8481: data <= 8'hFF;
            15'd8482: data <= 8'hFF;
            15'd8483: data <= 8'hFF;
            15'd8484: data <= 8'hFF;
            15'd8485: data <= 8'h80;
            15'd8486: data <= 8'h00;
            15'd8487: data <= 8'h00;
            15'd8488: data <= 8'h00;
            15'd8489: data <= 8'h00;
            15'd8490: data <= 8'h00;
            15'd8491: data <= 8'h00;
            15'd8492: data <= 8'h00;
            15'd8493: data <= 8'h00;
            15'd8494: data <= 8'h01;
            15'd8495: data <= 8'hFF;
            15'd8496: data <= 8'hFF;
            15'd8497: data <= 8'hFF;
            15'd8498: data <= 8'hFF;
            15'd8499: data <= 8'hFF;
            15'd8500: data <= 8'hFF;
            15'd8501: data <= 8'hFF;
            15'd8502: data <= 8'hFF;
            15'd8503: data <= 8'hFF;
            15'd8504: data <= 8'hFF;
            15'd8505: data <= 8'h8F;
            15'd8506: data <= 8'hFF;
            15'd8507: data <= 8'hFF;
            15'd8508: data <= 8'hFF;
            15'd8509: data <= 8'hFF;
            15'd8510: data <= 8'hFF;
            15'd8511: data <= 8'hFF;
            15'd8512: data <= 8'hFF;
            15'd8513: data <= 8'hFF;
            15'd8514: data <= 8'hFF;
            15'd8515: data <= 8'h80;
            15'd8516: data <= 8'h00;
            15'd8517: data <= 8'h00;
            15'd8518: data <= 8'h00;
            15'd8519: data <= 8'h00;
            15'd8520: data <= 8'h00;
            15'd8521: data <= 8'h00;
            15'd8522: data <= 8'h00;
            15'd8523: data <= 8'h00;
            15'd8524: data <= 8'h01;
            15'd8525: data <= 8'hFF;
            15'd8526: data <= 8'hFF;
            15'd8527: data <= 8'hFF;
            15'd8528: data <= 8'hFF;
            15'd8529: data <= 8'hFF;
            15'd8530: data <= 8'hFF;
            15'd8531: data <= 8'hFF;
            15'd8532: data <= 8'hFF;
            15'd8533: data <= 8'hFF;
            15'd8534: data <= 8'hFF;
            15'd8535: data <= 8'h1F;
            15'd8536: data <= 8'h7F;
            15'd8537: data <= 8'hFF;
            15'd8538: data <= 8'hFF;
            15'd8539: data <= 8'hFF;
            15'd8540: data <= 8'hFF;
            15'd8541: data <= 8'hFF;
            15'd8542: data <= 8'hFF;
            15'd8543: data <= 8'hFF;
            15'd8544: data <= 8'hFF;
            15'd8545: data <= 8'h80;
            15'd8546: data <= 8'h00;
            15'd8547: data <= 8'h00;
            15'd8548: data <= 8'h00;
            15'd8549: data <= 8'h00;
            15'd8550: data <= 8'h00;
            15'd8551: data <= 8'h00;
            15'd8552: data <= 8'h00;
            15'd8553: data <= 8'h00;
            15'd8554: data <= 8'h01;
            15'd8555: data <= 8'hFF;
            15'd8556: data <= 8'hFF;
            15'd8557: data <= 8'hFF;
            15'd8558: data <= 8'hFF;
            15'd8559: data <= 8'hFF;
            15'd8560: data <= 8'hFF;
            15'd8561: data <= 8'hFF;
            15'd8562: data <= 8'hFF;
            15'd8563: data <= 8'hFF;
            15'd8564: data <= 8'hFE;
            15'd8565: data <= 8'h1E;
            15'd8566: data <= 8'h3F;
            15'd8567: data <= 8'h9F;
            15'd8568: data <= 8'hFF;
            15'd8569: data <= 8'hFF;
            15'd8570: data <= 8'hFF;
            15'd8571: data <= 8'hFF;
            15'd8572: data <= 8'hFF;
            15'd8573: data <= 8'hFF;
            15'd8574: data <= 8'hFF;
            15'd8575: data <= 8'h80;
            15'd8576: data <= 8'h00;
            15'd8577: data <= 8'h00;
            15'd8578: data <= 8'h00;
            15'd8579: data <= 8'h00;
            15'd8580: data <= 8'h00;
            15'd8581: data <= 8'h00;
            15'd8582: data <= 8'h00;
            15'd8583: data <= 8'h00;
            15'd8584: data <= 8'h01;
            15'd8585: data <= 8'hFF;
            15'd8586: data <= 8'hFF;
            15'd8587: data <= 8'hFF;
            15'd8588: data <= 8'hFF;
            15'd8589: data <= 8'hFF;
            15'd8590: data <= 8'hFF;
            15'd8591: data <= 8'hFF;
            15'd8592: data <= 8'hFF;
            15'd8593: data <= 8'hFF;
            15'd8594: data <= 8'hFE;
            15'd8595: data <= 8'h3C;
            15'd8596: data <= 8'h7F;
            15'd8597: data <= 8'h1F;
            15'd8598: data <= 8'hFF;
            15'd8599: data <= 8'hFF;
            15'd8600: data <= 8'hFF;
            15'd8601: data <= 8'hFF;
            15'd8602: data <= 8'hFF;
            15'd8603: data <= 8'hFF;
            15'd8604: data <= 8'hFF;
            15'd8605: data <= 8'h80;
            15'd8606: data <= 8'h00;
            15'd8607: data <= 8'h00;
            15'd8608: data <= 8'h00;
            15'd8609: data <= 8'h00;
            15'd8610: data <= 8'h00;
            15'd8611: data <= 8'h00;
            15'd8612: data <= 8'h00;
            15'd8613: data <= 8'h00;
            15'd8614: data <= 8'h01;
            15'd8615: data <= 8'hFF;
            15'd8616: data <= 8'hFF;
            15'd8617: data <= 8'hFF;
            15'd8618: data <= 8'hFF;
            15'd8619: data <= 8'hFF;
            15'd8620: data <= 8'hFF;
            15'd8621: data <= 8'hFF;
            15'd8622: data <= 8'hFF;
            15'd8623: data <= 8'hFF;
            15'd8624: data <= 8'hFC;
            15'd8625: data <= 8'h7C;
            15'd8626: data <= 8'h7E;
            15'd8627: data <= 8'h1F;
            15'd8628: data <= 8'hFF;
            15'd8629: data <= 8'hFF;
            15'd8630: data <= 8'hFF;
            15'd8631: data <= 8'hFF;
            15'd8632: data <= 8'hFF;
            15'd8633: data <= 8'hFF;
            15'd8634: data <= 8'hFF;
            15'd8635: data <= 8'h80;
            15'd8636: data <= 8'h00;
            15'd8637: data <= 8'h00;
            15'd8638: data <= 8'h00;
            15'd8639: data <= 8'h00;
            15'd8640: data <= 8'h00;
            15'd8641: data <= 8'h00;
            15'd8642: data <= 8'h00;
            15'd8643: data <= 8'h00;
            15'd8644: data <= 8'h01;
            15'd8645: data <= 8'hFF;
            15'd8646: data <= 8'hFF;
            15'd8647: data <= 8'hFF;
            15'd8648: data <= 8'hFF;
            15'd8649: data <= 8'hFF;
            15'd8650: data <= 8'hFF;
            15'd8651: data <= 8'hFF;
            15'd8652: data <= 8'hFF;
            15'd8653: data <= 8'hFF;
            15'd8654: data <= 8'hFF;
            15'd8655: data <= 8'hF8;
            15'd8656: data <= 8'hFE;
            15'd8657: data <= 8'h3F;
            15'd8658: data <= 8'hFF;
            15'd8659: data <= 8'hFF;
            15'd8660: data <= 8'hFF;
            15'd8661: data <= 8'hFF;
            15'd8662: data <= 8'hFF;
            15'd8663: data <= 8'hFF;
            15'd8664: data <= 8'hFF;
            15'd8665: data <= 8'h80;
            15'd8666: data <= 8'h00;
            15'd8667: data <= 8'h00;
            15'd8668: data <= 8'h00;
            15'd8669: data <= 8'h00;
            15'd8670: data <= 8'h00;
            15'd8671: data <= 8'h00;
            15'd8672: data <= 8'h00;
            15'd8673: data <= 8'h00;
            15'd8674: data <= 8'h01;
            15'd8675: data <= 8'hFF;
            15'd8676: data <= 8'hFF;
            15'd8677: data <= 8'hFF;
            15'd8678: data <= 8'hFF;
            15'd8679: data <= 8'hFF;
            15'd8680: data <= 8'hFF;
            15'd8681: data <= 8'hFF;
            15'd8682: data <= 8'hFF;
            15'd8683: data <= 8'hFF;
            15'd8684: data <= 8'hFF;
            15'd8685: data <= 8'hF1;
            15'd8686: data <= 8'hFC;
            15'd8687: data <= 8'h7F;
            15'd8688: data <= 8'hFF;
            15'd8689: data <= 8'hFF;
            15'd8690: data <= 8'hFF;
            15'd8691: data <= 8'hFF;
            15'd8692: data <= 8'hFF;
            15'd8693: data <= 8'hFF;
            15'd8694: data <= 8'hFF;
            15'd8695: data <= 8'h80;
            15'd8696: data <= 8'h00;
            15'd8697: data <= 8'h00;
            15'd8698: data <= 8'h00;
            15'd8699: data <= 8'h00;
            15'd8700: data <= 8'h00;
            15'd8701: data <= 8'h00;
            15'd8702: data <= 8'h00;
            15'd8703: data <= 8'h00;
            15'd8704: data <= 8'h01;
            15'd8705: data <= 8'hFF;
            15'd8706: data <= 8'hFF;
            15'd8707: data <= 8'hFF;
            15'd8708: data <= 8'hFF;
            15'd8709: data <= 8'hFF;
            15'd8710: data <= 8'hFF;
            15'd8711: data <= 8'hFF;
            15'd8712: data <= 8'hFF;
            15'd8713: data <= 8'hFF;
            15'd8714: data <= 8'hFF;
            15'd8715: data <= 8'hF1;
            15'd8716: data <= 8'hF8;
            15'd8717: data <= 8'hFF;
            15'd8718: data <= 8'hFF;
            15'd8719: data <= 8'hFF;
            15'd8720: data <= 8'hFF;
            15'd8721: data <= 8'hFF;
            15'd8722: data <= 8'hFF;
            15'd8723: data <= 8'hFF;
            15'd8724: data <= 8'hFF;
            15'd8725: data <= 8'h80;
            15'd8726: data <= 8'h00;
            15'd8727: data <= 8'h00;
            15'd8728: data <= 8'h00;
            15'd8729: data <= 8'h00;
            15'd8730: data <= 8'h00;
            15'd8731: data <= 8'h00;
            15'd8732: data <= 8'h00;
            15'd8733: data <= 8'h00;
            15'd8734: data <= 8'h01;
            15'd8735: data <= 8'hFF;
            15'd8736: data <= 8'hFF;
            15'd8737: data <= 8'hFF;
            15'd8738: data <= 8'hFF;
            15'd8739: data <= 8'hFF;
            15'd8740: data <= 8'hFF;
            15'd8741: data <= 8'hFF;
            15'd8742: data <= 8'hFF;
            15'd8743: data <= 8'hFF;
            15'd8744: data <= 8'hFF;
            15'd8745: data <= 8'hE3;
            15'd8746: data <= 8'hF0;
            15'd8747: data <= 8'hFF;
            15'd8748: data <= 8'hFF;
            15'd8749: data <= 8'hFF;
            15'd8750: data <= 8'hFF;
            15'd8751: data <= 8'hFF;
            15'd8752: data <= 8'hFF;
            15'd8753: data <= 8'hFF;
            15'd8754: data <= 8'hFF;
            15'd8755: data <= 8'h80;
            15'd8756: data <= 8'h00;
            15'd8757: data <= 8'h00;
            15'd8758: data <= 8'h00;
            15'd8759: data <= 8'h00;
            15'd8760: data <= 8'h00;
            15'd8761: data <= 8'h00;
            15'd8762: data <= 8'h00;
            15'd8763: data <= 8'h00;
            15'd8764: data <= 8'h01;
            15'd8765: data <= 8'hFF;
            15'd8766: data <= 8'hFF;
            15'd8767: data <= 8'hFF;
            15'd8768: data <= 8'hFF;
            15'd8769: data <= 8'hFF;
            15'd8770: data <= 8'hFF;
            15'd8771: data <= 8'hFF;
            15'd8772: data <= 8'hFF;
            15'd8773: data <= 8'hFF;
            15'd8774: data <= 8'hFF;
            15'd8775: data <= 8'hE7;
            15'd8776: data <= 8'hF1;
            15'd8777: data <= 8'hFF;
            15'd8778: data <= 8'hFF;
            15'd8779: data <= 8'hFF;
            15'd8780: data <= 8'hFF;
            15'd8781: data <= 8'hFF;
            15'd8782: data <= 8'hFF;
            15'd8783: data <= 8'hFF;
            15'd8784: data <= 8'hFF;
            15'd8785: data <= 8'h80;
            15'd8786: data <= 8'h00;
            15'd8787: data <= 8'h00;
            15'd8788: data <= 8'h00;
            15'd8789: data <= 8'h00;
            15'd8790: data <= 8'h00;
            15'd8791: data <= 8'h00;
            15'd8792: data <= 8'h00;
            15'd8793: data <= 8'h00;
            15'd8794: data <= 8'h01;
            15'd8795: data <= 8'hFF;
            15'd8796: data <= 8'hFF;
            15'd8797: data <= 8'hFF;
            15'd8798: data <= 8'hFF;
            15'd8799: data <= 8'hFF;
            15'd8800: data <= 8'hFF;
            15'd8801: data <= 8'hFF;
            15'd8802: data <= 8'hFF;
            15'd8803: data <= 8'hC0;
            15'd8804: data <= 8'hFF;
            15'd8805: data <= 8'hEF;
            15'd8806: data <= 8'hE3;
            15'd8807: data <= 8'hFF;
            15'd8808: data <= 8'hFF;
            15'd8809: data <= 8'hFF;
            15'd8810: data <= 8'hFF;
            15'd8811: data <= 8'hFF;
            15'd8812: data <= 8'hFF;
            15'd8813: data <= 8'hFF;
            15'd8814: data <= 8'hFF;
            15'd8815: data <= 8'h80;
            15'd8816: data <= 8'h00;
            15'd8817: data <= 8'h00;
            15'd8818: data <= 8'h00;
            15'd8819: data <= 8'h00;
            15'd8820: data <= 8'h00;
            15'd8821: data <= 8'h00;
            15'd8822: data <= 8'h00;
            15'd8823: data <= 8'h00;
            15'd8824: data <= 8'h01;
            15'd8825: data <= 8'hFF;
            15'd8826: data <= 8'hFF;
            15'd8827: data <= 8'hFF;
            15'd8828: data <= 8'hFF;
            15'd8829: data <= 8'hFF;
            15'd8830: data <= 8'hFF;
            15'd8831: data <= 8'hFF;
            15'd8832: data <= 8'hE3;
            15'd8833: data <= 8'h80;
            15'd8834: data <= 8'h7F;
            15'd8835: data <= 8'hFF;
            15'd8836: data <= 8'hC3;
            15'd8837: data <= 8'hFF;
            15'd8838: data <= 8'hFF;
            15'd8839: data <= 8'hFF;
            15'd8840: data <= 8'hFF;
            15'd8841: data <= 8'hFF;
            15'd8842: data <= 8'hFF;
            15'd8843: data <= 8'hFF;
            15'd8844: data <= 8'hFF;
            15'd8845: data <= 8'h80;
            15'd8846: data <= 8'h00;
            15'd8847: data <= 8'h00;
            15'd8848: data <= 8'h00;
            15'd8849: data <= 8'h00;
            15'd8850: data <= 8'h00;
            15'd8851: data <= 8'h00;
            15'd8852: data <= 8'h00;
            15'd8853: data <= 8'h00;
            15'd8854: data <= 8'h01;
            15'd8855: data <= 8'hFF;
            15'd8856: data <= 8'hFF;
            15'd8857: data <= 8'hFF;
            15'd8858: data <= 8'hFF;
            15'd8859: data <= 8'hFF;
            15'd8860: data <= 8'hFF;
            15'd8861: data <= 8'hFF;
            15'd8862: data <= 8'h00;
            15'd8863: data <= 8'h00;
            15'd8864: data <= 8'h3F;
            15'd8865: data <= 8'hFF;
            15'd8866: data <= 8'hC7;
            15'd8867: data <= 8'hFF;
            15'd8868: data <= 8'hFF;
            15'd8869: data <= 8'hFF;
            15'd8870: data <= 8'hFF;
            15'd8871: data <= 8'hFF;
            15'd8872: data <= 8'hFF;
            15'd8873: data <= 8'hFF;
            15'd8874: data <= 8'hFF;
            15'd8875: data <= 8'h80;
            15'd8876: data <= 8'h00;
            15'd8877: data <= 8'h00;
            15'd8878: data <= 8'h00;
            15'd8879: data <= 8'h00;
            15'd8880: data <= 8'h00;
            15'd8881: data <= 8'h00;
            15'd8882: data <= 8'h00;
            15'd8883: data <= 8'h00;
            15'd8884: data <= 8'h01;
            15'd8885: data <= 8'hFF;
            15'd8886: data <= 8'hFF;
            15'd8887: data <= 8'hFF;
            15'd8888: data <= 8'hFF;
            15'd8889: data <= 8'hFF;
            15'd8890: data <= 8'hFF;
            15'd8891: data <= 8'hFF;
            15'd8892: data <= 8'h00;
            15'd8893: data <= 8'h04;
            15'd8894: data <= 8'h3F;
            15'd8895: data <= 8'hFF;
            15'd8896: data <= 8'h8F;
            15'd8897: data <= 8'hFF;
            15'd8898: data <= 8'hFF;
            15'd8899: data <= 8'hFF;
            15'd8900: data <= 8'hFF;
            15'd8901: data <= 8'hFF;
            15'd8902: data <= 8'hFF;
            15'd8903: data <= 8'hFF;
            15'd8904: data <= 8'hFF;
            15'd8905: data <= 8'h80;
            15'd8906: data <= 8'h00;
            15'd8907: data <= 8'h00;
            15'd8908: data <= 8'h00;
            15'd8909: data <= 8'h00;
            15'd8910: data <= 8'h00;
            15'd8911: data <= 8'h00;
            15'd8912: data <= 8'h00;
            15'd8913: data <= 8'h00;
            15'd8914: data <= 8'h01;
            15'd8915: data <= 8'hFF;
            15'd8916: data <= 8'hFF;
            15'd8917: data <= 8'hFF;
            15'd8918: data <= 8'hFF;
            15'd8919: data <= 8'hFF;
            15'd8920: data <= 8'hFF;
            15'd8921: data <= 8'hFE;
            15'd8922: data <= 8'h0C;
            15'd8923: data <= 8'h1E;
            15'd8924: data <= 8'h3F;
            15'd8925: data <= 8'hFF;
            15'd8926: data <= 8'h9F;
            15'd8927: data <= 8'hFF;
            15'd8928: data <= 8'hFF;
            15'd8929: data <= 8'hFF;
            15'd8930: data <= 8'hFF;
            15'd8931: data <= 8'hFF;
            15'd8932: data <= 8'hFF;
            15'd8933: data <= 8'hFF;
            15'd8934: data <= 8'hFF;
            15'd8935: data <= 8'h80;
            15'd8936: data <= 8'h00;
            15'd8937: data <= 8'h00;
            15'd8938: data <= 8'h00;
            15'd8939: data <= 8'h00;
            15'd8940: data <= 8'h00;
            15'd8941: data <= 8'h00;
            15'd8942: data <= 8'h00;
            15'd8943: data <= 8'h00;
            15'd8944: data <= 8'h01;
            15'd8945: data <= 8'hFF;
            15'd8946: data <= 8'hFF;
            15'd8947: data <= 8'hFF;
            15'd8948: data <= 8'hFF;
            15'd8949: data <= 8'hFF;
            15'd8950: data <= 8'hFF;
            15'd8951: data <= 8'hFE;
            15'd8952: data <= 8'h1E;
            15'd8953: data <= 8'h3E;
            15'd8954: data <= 8'h3F;
            15'd8955: data <= 8'hFF;
            15'd8956: data <= 8'h3F;
            15'd8957: data <= 8'hFF;
            15'd8958: data <= 8'hFF;
            15'd8959: data <= 8'hFF;
            15'd8960: data <= 8'hFF;
            15'd8961: data <= 8'hFF;
            15'd8962: data <= 8'hFF;
            15'd8963: data <= 8'hFF;
            15'd8964: data <= 8'hFF;
            15'd8965: data <= 8'h80;
            15'd8966: data <= 8'h00;
            15'd8967: data <= 8'h00;
            15'd8968: data <= 8'h00;
            15'd8969: data <= 8'h00;
            15'd8970: data <= 8'h00;
            15'd8971: data <= 8'h00;
            15'd8972: data <= 8'h00;
            15'd8973: data <= 8'h00;
            15'd8974: data <= 8'h01;
            15'd8975: data <= 8'hFF;
            15'd8976: data <= 8'hFF;
            15'd8977: data <= 8'hFF;
            15'd8978: data <= 8'hFF;
            15'd8979: data <= 8'hFF;
            15'd8980: data <= 8'hFF;
            15'd8981: data <= 8'hFE;
            15'd8982: data <= 8'h1F;
            15'd8983: data <= 8'hFE;
            15'd8984: data <= 8'h3F;
            15'd8985: data <= 8'hFF;
            15'd8986: data <= 8'h3F;
            15'd8987: data <= 8'hFF;
            15'd8988: data <= 8'hFF;
            15'd8989: data <= 8'hFF;
            15'd8990: data <= 8'hFF;
            15'd8991: data <= 8'hFF;
            15'd8992: data <= 8'hFF;
            15'd8993: data <= 8'hFF;
            15'd8994: data <= 8'hFF;
            15'd8995: data <= 8'h80;
            15'd8996: data <= 8'h00;
            15'd8997: data <= 8'h00;
            15'd8998: data <= 8'h00;
            15'd8999: data <= 8'h00;
            15'd9000: data <= 8'h00;
            15'd9001: data <= 8'h00;
            15'd9002: data <= 8'h00;
            15'd9003: data <= 8'h00;
            15'd9004: data <= 8'h01;
            15'd9005: data <= 8'hFF;
            15'd9006: data <= 8'hFF;
            15'd9007: data <= 8'hFF;
            15'd9008: data <= 8'hFF;
            15'd9009: data <= 8'hFF;
            15'd9010: data <= 8'hFF;
            15'd9011: data <= 8'hFE;
            15'd9012: data <= 8'h1F;
            15'd9013: data <= 8'hFC;
            15'd9014: data <= 8'h3F;
            15'd9015: data <= 8'hFE;
            15'd9016: data <= 8'h7F;
            15'd9017: data <= 8'hFF;
            15'd9018: data <= 8'hFF;
            15'd9019: data <= 8'hFF;
            15'd9020: data <= 8'hFF;
            15'd9021: data <= 8'hFF;
            15'd9022: data <= 8'hFF;
            15'd9023: data <= 8'hFF;
            15'd9024: data <= 8'hFF;
            15'd9025: data <= 8'h80;
            15'd9026: data <= 8'h00;
            15'd9027: data <= 8'h00;
            15'd9028: data <= 8'h00;
            15'd9029: data <= 8'h00;
            15'd9030: data <= 8'h00;
            15'd9031: data <= 8'h00;
            15'd9032: data <= 8'h00;
            15'd9033: data <= 8'h00;
            15'd9034: data <= 8'h01;
            15'd9035: data <= 8'hFF;
            15'd9036: data <= 8'hFF;
            15'd9037: data <= 8'hFF;
            15'd9038: data <= 8'hFF;
            15'd9039: data <= 8'hFF;
            15'd9040: data <= 8'hFF;
            15'd9041: data <= 8'hFE;
            15'd9042: data <= 8'h1F;
            15'd9043: data <= 8'hFC;
            15'd9044: data <= 8'h3F;
            15'd9045: data <= 8'hFC;
            15'd9046: data <= 8'hFF;
            15'd9047: data <= 8'hFF;
            15'd9048: data <= 8'hFF;
            15'd9049: data <= 8'hFF;
            15'd9050: data <= 8'hFF;
            15'd9051: data <= 8'hFF;
            15'd9052: data <= 8'hFF;
            15'd9053: data <= 8'hFF;
            15'd9054: data <= 8'hFF;
            15'd9055: data <= 8'h80;
            15'd9056: data <= 8'h00;
            15'd9057: data <= 8'h00;
            15'd9058: data <= 8'h00;
            15'd9059: data <= 8'h00;
            15'd9060: data <= 8'h00;
            15'd9061: data <= 8'h00;
            15'd9062: data <= 8'h00;
            15'd9063: data <= 8'h00;
            15'd9064: data <= 8'h01;
            15'd9065: data <= 8'hFF;
            15'd9066: data <= 8'hFF;
            15'd9067: data <= 8'hFF;
            15'd9068: data <= 8'hFF;
            15'd9069: data <= 8'hFF;
            15'd9070: data <= 8'hFF;
            15'd9071: data <= 8'hFF;
            15'd9072: data <= 8'h0F;
            15'd9073: data <= 8'hF8;
            15'd9074: data <= 8'h7F;
            15'd9075: data <= 8'hFD;
            15'd9076: data <= 8'hFF;
            15'd9077: data <= 8'hFF;
            15'd9078: data <= 8'hFF;
            15'd9079: data <= 8'hFF;
            15'd9080: data <= 8'hFF;
            15'd9081: data <= 8'hFF;
            15'd9082: data <= 8'hFF;
            15'd9083: data <= 8'hFF;
            15'd9084: data <= 8'hFF;
            15'd9085: data <= 8'h80;
            15'd9086: data <= 8'h00;
            15'd9087: data <= 8'h00;
            15'd9088: data <= 8'h00;
            15'd9089: data <= 8'h00;
            15'd9090: data <= 8'h00;
            15'd9091: data <= 8'h00;
            15'd9092: data <= 8'h00;
            15'd9093: data <= 8'h00;
            15'd9094: data <= 8'h01;
            15'd9095: data <= 8'hFF;
            15'd9096: data <= 8'hFF;
            15'd9097: data <= 8'hFF;
            15'd9098: data <= 8'hFF;
            15'd9099: data <= 8'hFF;
            15'd9100: data <= 8'hFF;
            15'd9101: data <= 8'hFF;
            15'd9102: data <= 8'h87;
            15'd9103: data <= 8'hF8;
            15'd9104: data <= 8'h7F;
            15'd9105: data <= 8'hF9;
            15'd9106: data <= 8'hFF;
            15'd9107: data <= 8'hFF;
            15'd9108: data <= 8'hFF;
            15'd9109: data <= 8'hFF;
            15'd9110: data <= 8'hFF;
            15'd9111: data <= 8'hFF;
            15'd9112: data <= 8'hFF;
            15'd9113: data <= 8'hFF;
            15'd9114: data <= 8'hFF;
            15'd9115: data <= 8'h80;
            15'd9116: data <= 8'h00;
            15'd9117: data <= 8'h00;
            15'd9118: data <= 8'h00;
            15'd9119: data <= 8'h00;
            15'd9120: data <= 8'h00;
            15'd9121: data <= 8'h00;
            15'd9122: data <= 8'h00;
            15'd9123: data <= 8'h00;
            15'd9124: data <= 8'h01;
            15'd9125: data <= 8'hFF;
            15'd9126: data <= 8'hFF;
            15'd9127: data <= 8'hFF;
            15'd9128: data <= 8'hFF;
            15'd9129: data <= 8'hFF;
            15'd9130: data <= 8'hFF;
            15'd9131: data <= 8'hFF;
            15'd9132: data <= 8'h83;
            15'd9133: data <= 8'hF0;
            15'd9134: data <= 8'hFF;
            15'd9135: data <= 8'hFF;
            15'd9136: data <= 8'hFF;
            15'd9137: data <= 8'hFF;
            15'd9138: data <= 8'hFF;
            15'd9139: data <= 8'hFF;
            15'd9140: data <= 8'hFF;
            15'd9141: data <= 8'hFF;
            15'd9142: data <= 8'hFF;
            15'd9143: data <= 8'hFF;
            15'd9144: data <= 8'hFF;
            15'd9145: data <= 8'h80;
            15'd9146: data <= 8'h00;
            15'd9147: data <= 8'h00;
            15'd9148: data <= 8'h00;
            15'd9149: data <= 8'h00;
            15'd9150: data <= 8'h00;
            15'd9151: data <= 8'h00;
            15'd9152: data <= 8'h00;
            15'd9153: data <= 8'h00;
            15'd9154: data <= 8'h01;
            15'd9155: data <= 8'hFF;
            15'd9156: data <= 8'hFF;
            15'd9157: data <= 8'hFF;
            15'd9158: data <= 8'hFF;
            15'd9159: data <= 8'hFF;
            15'd9160: data <= 8'hFF;
            15'd9161: data <= 8'hFF;
            15'd9162: data <= 8'hC1;
            15'd9163: data <= 8'hE0;
            15'd9164: data <= 8'hFF;
            15'd9165: data <= 8'hFF;
            15'd9166: data <= 8'hFF;
            15'd9167: data <= 8'hFF;
            15'd9168: data <= 8'hFF;
            15'd9169: data <= 8'hFF;
            15'd9170: data <= 8'hFF;
            15'd9171: data <= 8'hFF;
            15'd9172: data <= 8'hFF;
            15'd9173: data <= 8'hFF;
            15'd9174: data <= 8'hFF;
            15'd9175: data <= 8'h80;
            15'd9176: data <= 8'h00;
            15'd9177: data <= 8'h00;
            15'd9178: data <= 8'h00;
            15'd9179: data <= 8'h00;
            15'd9180: data <= 8'h00;
            15'd9181: data <= 8'h00;
            15'd9182: data <= 8'h00;
            15'd9183: data <= 8'h00;
            15'd9184: data <= 8'h01;
            15'd9185: data <= 8'hFF;
            15'd9186: data <= 8'hFF;
            15'd9187: data <= 8'hFF;
            15'd9188: data <= 8'hFF;
            15'd9189: data <= 8'hFF;
            15'd9190: data <= 8'hFF;
            15'd9191: data <= 8'hFF;
            15'd9192: data <= 8'hE0;
            15'd9193: data <= 8'h41;
            15'd9194: data <= 8'hFF;
            15'd9195: data <= 8'hFF;
            15'd9196: data <= 8'hFF;
            15'd9197: data <= 8'hFF;
            15'd9198: data <= 8'hFF;
            15'd9199: data <= 8'hFF;
            15'd9200: data <= 8'hFF;
            15'd9201: data <= 8'hFF;
            15'd9202: data <= 8'hFF;
            15'd9203: data <= 8'hFF;
            15'd9204: data <= 8'hFF;
            15'd9205: data <= 8'h80;
            15'd9206: data <= 8'h00;
            15'd9207: data <= 8'h00;
            15'd9208: data <= 8'h00;
            15'd9209: data <= 8'h00;
            15'd9210: data <= 8'h00;
            15'd9211: data <= 8'h00;
            15'd9212: data <= 8'h00;
            15'd9213: data <= 8'h00;
            15'd9214: data <= 8'h01;
            15'd9215: data <= 8'hFF;
            15'd9216: data <= 8'hFF;
            15'd9217: data <= 8'hFF;
            15'd9218: data <= 8'hFF;
            15'd9219: data <= 8'hFF;
            15'd9220: data <= 8'hFF;
            15'd9221: data <= 8'hFF;
            15'd9222: data <= 8'hF8;
            15'd9223: data <= 8'h03;
            15'd9224: data <= 8'hFF;
            15'd9225: data <= 8'hFF;
            15'd9226: data <= 8'hFF;
            15'd9227: data <= 8'hFF;
            15'd9228: data <= 8'hFF;
            15'd9229: data <= 8'hFF;
            15'd9230: data <= 8'hFF;
            15'd9231: data <= 8'hFF;
            15'd9232: data <= 8'hFF;
            15'd9233: data <= 8'hFF;
            15'd9234: data <= 8'hFF;
            15'd9235: data <= 8'h80;
            15'd9236: data <= 8'h00;
            15'd9237: data <= 8'h00;
            15'd9238: data <= 8'h00;
            15'd9239: data <= 8'h00;
            15'd9240: data <= 8'h00;
            15'd9241: data <= 8'h00;
            15'd9242: data <= 8'h00;
            15'd9243: data <= 8'h00;
            15'd9244: data <= 8'h01;
            15'd9245: data <= 8'hFF;
            15'd9246: data <= 8'hFF;
            15'd9247: data <= 8'hFF;
            15'd9248: data <= 8'hFF;
            15'd9249: data <= 8'hFF;
            15'd9250: data <= 8'hFF;
            15'd9251: data <= 8'hFF;
            15'd9252: data <= 8'hEC;
            15'd9253: data <= 8'h07;
            15'd9254: data <= 8'hFF;
            15'd9255: data <= 8'hFF;
            15'd9256: data <= 8'hFF;
            15'd9257: data <= 8'hFF;
            15'd9258: data <= 8'hFF;
            15'd9259: data <= 8'hFF;
            15'd9260: data <= 8'hFF;
            15'd9261: data <= 8'hFF;
            15'd9262: data <= 8'hFF;
            15'd9263: data <= 8'hFF;
            15'd9264: data <= 8'hFF;
            15'd9265: data <= 8'h80;
            15'd9266: data <= 8'h00;
            15'd9267: data <= 8'h00;
            15'd9268: data <= 8'h00;
            15'd9269: data <= 8'h00;
            15'd9270: data <= 8'h00;
            15'd9271: data <= 8'h00;
            15'd9272: data <= 8'h00;
            15'd9273: data <= 8'h00;
            15'd9274: data <= 8'h01;
            15'd9275: data <= 8'hFF;
            15'd9276: data <= 8'hFF;
            15'd9277: data <= 8'hFF;
            15'd9278: data <= 8'hFF;
            15'd9279: data <= 8'hFF;
            15'd9280: data <= 8'hFF;
            15'd9281: data <= 8'hFF;
            15'd9282: data <= 8'hF6;
            15'd9283: data <= 8'h0F;
            15'd9284: data <= 8'hFF;
            15'd9285: data <= 8'hFF;
            15'd9286: data <= 8'hFF;
            15'd9287: data <= 8'hFF;
            15'd9288: data <= 8'hFF;
            15'd9289: data <= 8'hFF;
            15'd9290: data <= 8'hFF;
            15'd9291: data <= 8'hFF;
            15'd9292: data <= 8'hFF;
            15'd9293: data <= 8'hFF;
            15'd9294: data <= 8'hFF;
            15'd9295: data <= 8'h80;
            15'd9296: data <= 8'h00;
            15'd9297: data <= 8'h00;
            15'd9298: data <= 8'h00;
            15'd9299: data <= 8'h00;
            15'd9300: data <= 8'h00;
            15'd9301: data <= 8'h00;
            15'd9302: data <= 8'h00;
            15'd9303: data <= 8'h00;
            15'd9304: data <= 8'h01;
            15'd9305: data <= 8'hFF;
            15'd9306: data <= 8'hFD;
            15'd9307: data <= 8'hFF;
            15'd9308: data <= 8'hFF;
            15'd9309: data <= 8'hFF;
            15'd9310: data <= 8'hFF;
            15'd9311: data <= 8'hFF;
            15'd9312: data <= 8'hFF;
            15'd9313: data <= 8'hFF;
            15'd9314: data <= 8'hFF;
            15'd9315: data <= 8'hFF;
            15'd9316: data <= 8'hFF;
            15'd9317: data <= 8'hFF;
            15'd9318: data <= 8'hFF;
            15'd9319: data <= 8'hFF;
            15'd9320: data <= 8'hFF;
            15'd9321: data <= 8'hFF;
            15'd9322: data <= 8'hFF;
            15'd9323: data <= 8'hFF;
            15'd9324: data <= 8'hFF;
            15'd9325: data <= 8'h80;
            15'd9326: data <= 8'h00;
            15'd9327: data <= 8'h00;
            15'd9328: data <= 8'h00;
            15'd9329: data <= 8'h00;
            15'd9330: data <= 8'h00;
            15'd9331: data <= 8'h00;
            15'd9332: data <= 8'h00;
            15'd9333: data <= 8'h00;
            15'd9334: data <= 8'h01;
            15'd9335: data <= 8'hFF;
            15'd9336: data <= 8'hFF;
            15'd9337: data <= 8'hFF;
            15'd9338: data <= 8'hFF;
            15'd9339: data <= 8'hFF;
            15'd9340: data <= 8'hFF;
            15'd9341: data <= 8'hFF;
            15'd9342: data <= 8'hFF;
            15'd9343: data <= 8'hFF;
            15'd9344: data <= 8'hFF;
            15'd9345: data <= 8'hFF;
            15'd9346: data <= 8'hFF;
            15'd9347: data <= 8'hFF;
            15'd9348: data <= 8'hFF;
            15'd9349: data <= 8'hFF;
            15'd9350: data <= 8'hFF;
            15'd9351: data <= 8'hFF;
            15'd9352: data <= 8'hFF;
            15'd9353: data <= 8'hFF;
            15'd9354: data <= 8'hFF;
            15'd9355: data <= 8'h80;
            15'd9356: data <= 8'h00;
            15'd9357: data <= 8'h00;
            15'd9358: data <= 8'h00;
            15'd9359: data <= 8'h00;
            15'd9360: data <= 8'h00;
            15'd9361: data <= 8'h00;
            15'd9362: data <= 8'h00;
            15'd9363: data <= 8'h00;
            15'd9364: data <= 8'h01;
            15'd9365: data <= 8'hFF;
            15'd9366: data <= 8'hFF;
            15'd9367: data <= 8'hFF;
            15'd9368: data <= 8'hFF;
            15'd9369: data <= 8'hFF;
            15'd9370: data <= 8'hFF;
            15'd9371: data <= 8'hFF;
            15'd9372: data <= 8'hFF;
            15'd9373: data <= 8'hFF;
            15'd9374: data <= 8'hFF;
            15'd9375: data <= 8'hFF;
            15'd9376: data <= 8'hFF;
            15'd9377: data <= 8'hFF;
            15'd9378: data <= 8'hFF;
            15'd9379: data <= 8'hFF;
            15'd9380: data <= 8'hFF;
            15'd9381: data <= 8'hFF;
            15'd9382: data <= 8'hFF;
            15'd9383: data <= 8'hFF;
            15'd9384: data <= 8'hFF;
            15'd9385: data <= 8'h80;
            15'd9386: data <= 8'h00;
            15'd9387: data <= 8'h00;
            15'd9388: data <= 8'h00;
            15'd9389: data <= 8'h00;
            15'd9390: data <= 8'h00;
            15'd9391: data <= 8'h00;
            15'd9392: data <= 8'h00;
            15'd9393: data <= 8'h00;
            15'd9394: data <= 8'h01;
            15'd9395: data <= 8'hFF;
            15'd9396: data <= 8'hFF;
            15'd9397: data <= 8'hFF;
            15'd9398: data <= 8'hFF;
            15'd9399: data <= 8'hFF;
            15'd9400: data <= 8'hFF;
            15'd9401: data <= 8'hFF;
            15'd9402: data <= 8'hFF;
            15'd9403: data <= 8'hFF;
            15'd9404: data <= 8'hFF;
            15'd9405: data <= 8'hFF;
            15'd9406: data <= 8'hFF;
            15'd9407: data <= 8'hFF;
            15'd9408: data <= 8'hFF;
            15'd9409: data <= 8'hFF;
            15'd9410: data <= 8'hFF;
            15'd9411: data <= 8'hFF;
            15'd9412: data <= 8'hFF;
            15'd9413: data <= 8'hFF;
            15'd9414: data <= 8'hFF;
            15'd9415: data <= 8'h80;
            15'd9416: data <= 8'h00;
            15'd9417: data <= 8'h00;
            15'd9418: data <= 8'h00;
            15'd9419: data <= 8'h00;
            15'd9420: data <= 8'h00;
            15'd9421: data <= 8'h00;
            15'd9422: data <= 8'h00;
            15'd9423: data <= 8'h00;
            15'd9424: data <= 8'h01;
            15'd9425: data <= 8'hFF;
            15'd9426: data <= 8'hFF;
            15'd9427: data <= 8'hFF;
            15'd9428: data <= 8'hFF;
            15'd9429: data <= 8'hFF;
            15'd9430: data <= 8'hFF;
            15'd9431: data <= 8'hFF;
            15'd9432: data <= 8'hFF;
            15'd9433: data <= 8'hFF;
            15'd9434: data <= 8'hFF;
            15'd9435: data <= 8'hFF;
            15'd9436: data <= 8'hFF;
            15'd9437: data <= 8'hFF;
            15'd9438: data <= 8'hFF;
            15'd9439: data <= 8'hFF;
            15'd9440: data <= 8'hFF;
            15'd9441: data <= 8'hFF;
            15'd9442: data <= 8'hFF;
            15'd9443: data <= 8'hFF;
            15'd9444: data <= 8'hFF;
            15'd9445: data <= 8'h80;
            15'd9446: data <= 8'h00;
            15'd9447: data <= 8'h00;
            15'd9448: data <= 8'h00;
            15'd9449: data <= 8'h00;
            15'd9450: data <= 8'h00;
            15'd9451: data <= 8'h00;
            15'd9452: data <= 8'h00;
            15'd9453: data <= 8'h00;
            15'd9454: data <= 8'h01;
            15'd9455: data <= 8'hFF;
            15'd9456: data <= 8'hFF;
            15'd9457: data <= 8'hFF;
            15'd9458: data <= 8'hFF;
            15'd9459: data <= 8'hFF;
            15'd9460: data <= 8'hFF;
            15'd9461: data <= 8'hFF;
            15'd9462: data <= 8'hFF;
            15'd9463: data <= 8'hFF;
            15'd9464: data <= 8'hFF;
            15'd9465: data <= 8'hFF;
            15'd9466: data <= 8'hFF;
            15'd9467: data <= 8'hFF;
            15'd9468: data <= 8'hFF;
            15'd9469: data <= 8'hFF;
            15'd9470: data <= 8'hFF;
            15'd9471: data <= 8'hFF;
            15'd9472: data <= 8'hFF;
            15'd9473: data <= 8'hFF;
            15'd9474: data <= 8'hFF;
            15'd9475: data <= 8'h80;
            15'd9476: data <= 8'h00;
            15'd9477: data <= 8'h00;
            15'd9478: data <= 8'h00;
            15'd9479: data <= 8'h00;
            15'd9480: data <= 8'h00;
            15'd9481: data <= 8'h00;
            15'd9482: data <= 8'h00;
            15'd9483: data <= 8'h00;
            15'd9484: data <= 8'h01;
            15'd9485: data <= 8'hFF;
            15'd9486: data <= 8'hFF;
            15'd9487: data <= 8'hFF;
            15'd9488: data <= 8'hFF;
            15'd9489: data <= 8'hFF;
            15'd9490: data <= 8'hFF;
            15'd9491: data <= 8'hFF;
            15'd9492: data <= 8'hFF;
            15'd9493: data <= 8'hFF;
            15'd9494: data <= 8'hFF;
            15'd9495: data <= 8'hFF;
            15'd9496: data <= 8'hFF;
            15'd9497: data <= 8'hFF;
            15'd9498: data <= 8'hFF;
            15'd9499: data <= 8'hFF;
            15'd9500: data <= 8'hFF;
            15'd9501: data <= 8'hFF;
            15'd9502: data <= 8'hFF;
            15'd9503: data <= 8'hFF;
            15'd9504: data <= 8'hFF;
            15'd9505: data <= 8'h80;
            15'd9506: data <= 8'h00;
            15'd9507: data <= 8'h00;
            15'd9508: data <= 8'h00;
            15'd9509: data <= 8'h00;
            15'd9510: data <= 8'h00;
            15'd9511: data <= 8'h00;
            15'd9512: data <= 8'h00;
            15'd9513: data <= 8'h00;
            15'd9514: data <= 8'h01;
            15'd9515: data <= 8'hFF;
            15'd9516: data <= 8'hFF;
            15'd9517: data <= 8'hFF;
            15'd9518: data <= 8'hFF;
            15'd9519: data <= 8'hFF;
            15'd9520: data <= 8'hFF;
            15'd9521: data <= 8'hFF;
            15'd9522: data <= 8'hFF;
            15'd9523: data <= 8'hFF;
            15'd9524: data <= 8'hFF;
            15'd9525: data <= 8'hFF;
            15'd9526: data <= 8'hFF;
            15'd9527: data <= 8'hFF;
            15'd9528: data <= 8'hFF;
            15'd9529: data <= 8'hFF;
            15'd9530: data <= 8'hFF;
            15'd9531: data <= 8'hFF;
            15'd9532: data <= 8'hFF;
            15'd9533: data <= 8'hFF;
            15'd9534: data <= 8'hFF;
            15'd9535: data <= 8'h80;
            15'd9536: data <= 8'h00;
            15'd9537: data <= 8'h00;
            15'd9538: data <= 8'h00;
            15'd9539: data <= 8'h00;
            15'd9540: data <= 8'h00;
            15'd9541: data <= 8'h00;
            15'd9542: data <= 8'h00;
            15'd9543: data <= 8'h00;
            15'd9544: data <= 8'h01;
            15'd9545: data <= 8'hFF;
            15'd9546: data <= 8'hFF;
            15'd9547: data <= 8'hFF;
            15'd9548: data <= 8'hFF;
            15'd9549: data <= 8'hFF;
            15'd9550: data <= 8'hFF;
            15'd9551: data <= 8'hFF;
            15'd9552: data <= 8'hFF;
            15'd9553: data <= 8'hFF;
            15'd9554: data <= 8'hFF;
            15'd9555: data <= 8'hFF;
            15'd9556: data <= 8'hFF;
            15'd9557: data <= 8'hFF;
            15'd9558: data <= 8'hFF;
            15'd9559: data <= 8'hFF;
            15'd9560: data <= 8'hFF;
            15'd9561: data <= 8'hFF;
            15'd9562: data <= 8'hFF;
            15'd9563: data <= 8'hFF;
            15'd9564: data <= 8'hFF;
            15'd9565: data <= 8'h80;
            15'd9566: data <= 8'h00;
            15'd9567: data <= 8'h00;
            15'd9568: data <= 8'h00;
            15'd9569: data <= 8'h00;
            15'd9570: data <= 8'h00;
            15'd9571: data <= 8'h00;
            15'd9572: data <= 8'h00;
            15'd9573: data <= 8'h00;
            15'd9574: data <= 8'h01;
            15'd9575: data <= 8'hFF;
            15'd9576: data <= 8'hFF;
            15'd9577: data <= 8'hFF;
            15'd9578: data <= 8'hFF;
            15'd9579: data <= 8'hFF;
            15'd9580: data <= 8'hFF;
            15'd9581: data <= 8'hFF;
            15'd9582: data <= 8'hFF;
            15'd9583: data <= 8'hFF;
            15'd9584: data <= 8'hFF;
            15'd9585: data <= 8'hFF;
            15'd9586: data <= 8'hFF;
            15'd9587: data <= 8'hFF;
            15'd9588: data <= 8'hFF;
            15'd9589: data <= 8'hFF;
            15'd9590: data <= 8'hFF;
            15'd9591: data <= 8'hFF;
            15'd9592: data <= 8'hFF;
            15'd9593: data <= 8'hFF;
            15'd9594: data <= 8'hFF;
            15'd9595: data <= 8'h80;
            15'd9596: data <= 8'h00;
            15'd9597: data <= 8'h00;
            15'd9598: data <= 8'h00;
            15'd9599: data <= 8'h00;
            15'd9600: data <= 8'h00;
            15'd9601: data <= 8'h00;
            15'd9602: data <= 8'h00;
            15'd9603: data <= 8'h00;
            15'd9604: data <= 8'h01;
            15'd9605: data <= 8'hFF;
            15'd9606: data <= 8'hFF;
            15'd9607: data <= 8'hFF;
            15'd9608: data <= 8'hFF;
            15'd9609: data <= 8'hFF;
            15'd9610: data <= 8'hFF;
            15'd9611: data <= 8'hFF;
            15'd9612: data <= 8'hFF;
            15'd9613: data <= 8'hFF;
            15'd9614: data <= 8'hFF;
            15'd9615: data <= 8'hFF;
            15'd9616: data <= 8'hFF;
            15'd9617: data <= 8'hFF;
            15'd9618: data <= 8'hFF;
            15'd9619: data <= 8'hFF;
            15'd9620: data <= 8'hFF;
            15'd9621: data <= 8'hFF;
            15'd9622: data <= 8'hFF;
            15'd9623: data <= 8'hFF;
            15'd9624: data <= 8'hFF;
            15'd9625: data <= 8'h80;
            15'd9626: data <= 8'h00;
            15'd9627: data <= 8'h00;
            15'd9628: data <= 8'h00;
            15'd9629: data <= 8'h00;
            15'd9630: data <= 8'h00;
            15'd9631: data <= 8'h00;
            15'd9632: data <= 8'h00;
            15'd9633: data <= 8'h00;
            15'd9634: data <= 8'h01;
            15'd9635: data <= 8'hFF;
            15'd9636: data <= 8'hFF;
            15'd9637: data <= 8'hFF;
            15'd9638: data <= 8'hFF;
            15'd9639: data <= 8'hFF;
            15'd9640: data <= 8'hFF;
            15'd9641: data <= 8'hFF;
            15'd9642: data <= 8'hFF;
            15'd9643: data <= 8'hFF;
            15'd9644: data <= 8'hFF;
            15'd9645: data <= 8'hFF;
            15'd9646: data <= 8'hFF;
            15'd9647: data <= 8'hFF;
            15'd9648: data <= 8'hFF;
            15'd9649: data <= 8'hFF;
            15'd9650: data <= 8'hFF;
            15'd9651: data <= 8'hFF;
            15'd9652: data <= 8'hFF;
            15'd9653: data <= 8'hFF;
            15'd9654: data <= 8'hFF;
            15'd9655: data <= 8'h80;
            15'd9656: data <= 8'h00;
            15'd9657: data <= 8'h00;
            15'd9658: data <= 8'h00;
            15'd9659: data <= 8'h00;
            15'd9660: data <= 8'h00;
            15'd9661: data <= 8'h00;
            15'd9662: data <= 8'h00;
            15'd9663: data <= 8'h00;
            15'd9664: data <= 8'h01;
            15'd9665: data <= 8'hFF;
            15'd9666: data <= 8'hFF;
            15'd9667: data <= 8'hFF;
            15'd9668: data <= 8'hFF;
            15'd9669: data <= 8'hFF;
            15'd9670: data <= 8'hFF;
            15'd9671: data <= 8'hFF;
            15'd9672: data <= 8'hFF;
            15'd9673: data <= 8'hFF;
            15'd9674: data <= 8'hFF;
            15'd9675: data <= 8'hFF;
            15'd9676: data <= 8'hFF;
            15'd9677: data <= 8'hFF;
            15'd9678: data <= 8'hFF;
            15'd9679: data <= 8'hFF;
            15'd9680: data <= 8'hFF;
            15'd9681: data <= 8'hFF;
            15'd9682: data <= 8'hFF;
            15'd9683: data <= 8'hFF;
            15'd9684: data <= 8'hFF;
            15'd9685: data <= 8'h80;
            15'd9686: data <= 8'h00;
            15'd9687: data <= 8'h00;
            15'd9688: data <= 8'h00;
            15'd9689: data <= 8'h00;
            15'd9690: data <= 8'h00;
            15'd9691: data <= 8'h00;
            15'd9692: data <= 8'h00;
            15'd9693: data <= 8'h00;
            15'd9694: data <= 8'h01;
            15'd9695: data <= 8'hFF;
            15'd9696: data <= 8'hFF;
            15'd9697: data <= 8'hFF;
            15'd9698: data <= 8'hFF;
            15'd9699: data <= 8'hFF;
            15'd9700: data <= 8'hFF;
            15'd9701: data <= 8'hFF;
            15'd9702: data <= 8'hFF;
            15'd9703: data <= 8'hFF;
            15'd9704: data <= 8'hFF;
            15'd9705: data <= 8'hFF;
            15'd9706: data <= 8'hFF;
            15'd9707: data <= 8'hFF;
            15'd9708: data <= 8'hFF;
            15'd9709: data <= 8'hFF;
            15'd9710: data <= 8'hFF;
            15'd9711: data <= 8'hFF;
            15'd9712: data <= 8'hFF;
            15'd9713: data <= 8'hFF;
            15'd9714: data <= 8'hFF;
            15'd9715: data <= 8'h80;
            15'd9716: data <= 8'h00;
            15'd9717: data <= 8'h00;
            15'd9718: data <= 8'h00;
            15'd9719: data <= 8'h00;
            15'd9720: data <= 8'h00;
            15'd9721: data <= 8'h00;
            15'd9722: data <= 8'h00;
            15'd9723: data <= 8'h00;
            15'd9724: data <= 8'h01;
            15'd9725: data <= 8'hFF;
            15'd9726: data <= 8'hFF;
            15'd9727: data <= 8'hFF;
            15'd9728: data <= 8'hFF;
            15'd9729: data <= 8'hFF;
            15'd9730: data <= 8'hFF;
            15'd9731: data <= 8'hFF;
            15'd9732: data <= 8'hFF;
            15'd9733: data <= 8'hEF;
            15'd9734: data <= 8'hFF;
            15'd9735: data <= 8'hF3;
            15'd9736: data <= 8'hFF;
            15'd9737: data <= 8'hFF;
            15'd9738: data <= 8'hFF;
            15'd9739: data <= 8'hFF;
            15'd9740: data <= 8'hFF;
            15'd9741: data <= 8'hFF;
            15'd9742: data <= 8'hFF;
            15'd9743: data <= 8'hFF;
            15'd9744: data <= 8'hFF;
            15'd9745: data <= 8'h80;
            15'd9746: data <= 8'h00;
            15'd9747: data <= 8'h00;
            15'd9748: data <= 8'h00;
            15'd9749: data <= 8'h00;
            15'd9750: data <= 8'h00;
            15'd9751: data <= 8'h00;
            15'd9752: data <= 8'h00;
            15'd9753: data <= 8'h00;
            15'd9754: data <= 8'h01;
            15'd9755: data <= 8'hFF;
            15'd9756: data <= 8'hFF;
            15'd9757: data <= 8'hFF;
            15'd9758: data <= 8'hFF;
            15'd9759: data <= 8'hFF;
            15'd9760: data <= 8'hFF;
            15'd9761: data <= 8'hFF;
            15'd9762: data <= 8'hFC;
            15'd9763: data <= 8'hC7;
            15'd9764: data <= 8'hFF;
            15'd9765: data <= 8'hF0;
            15'd9766: data <= 8'h03;
            15'd9767: data <= 8'hFF;
            15'd9768: data <= 8'hFF;
            15'd9769: data <= 8'hFF;
            15'd9770: data <= 8'hFF;
            15'd9771: data <= 8'hFF;
            15'd9772: data <= 8'hFF;
            15'd9773: data <= 8'hFF;
            15'd9774: data <= 8'hFF;
            15'd9775: data <= 8'h80;
            15'd9776: data <= 8'h00;
            15'd9777: data <= 8'h00;
            15'd9778: data <= 8'h00;
            15'd9779: data <= 8'h00;
            15'd9780: data <= 8'h00;
            15'd9781: data <= 8'h00;
            15'd9782: data <= 8'h00;
            15'd9783: data <= 8'h00;
            15'd9784: data <= 8'h01;
            15'd9785: data <= 8'hFF;
            15'd9786: data <= 8'hFF;
            15'd9787: data <= 8'hFF;
            15'd9788: data <= 8'hFF;
            15'd9789: data <= 8'hFF;
            15'd9790: data <= 8'hFF;
            15'd9791: data <= 8'hFF;
            15'd9792: data <= 8'hFC;
            15'd9793: data <= 8'h47;
            15'd9794: data <= 8'hFF;
            15'd9795: data <= 8'hE0;
            15'd9796: data <= 8'h01;
            15'd9797: data <= 8'hFF;
            15'd9798: data <= 8'hFF;
            15'd9799: data <= 8'hFF;
            15'd9800: data <= 8'hFF;
            15'd9801: data <= 8'hFF;
            15'd9802: data <= 8'hFF;
            15'd9803: data <= 8'hFF;
            15'd9804: data <= 8'hFF;
            15'd9805: data <= 8'h80;
            15'd9806: data <= 8'h00;
            15'd9807: data <= 8'h00;
            15'd9808: data <= 8'h00;
            15'd9809: data <= 8'h00;
            15'd9810: data <= 8'h00;
            15'd9811: data <= 8'h00;
            15'd9812: data <= 8'h00;
            15'd9813: data <= 8'h00;
            15'd9814: data <= 8'h01;
            15'd9815: data <= 8'hFF;
            15'd9816: data <= 8'hFF;
            15'd9817: data <= 8'hFF;
            15'd9818: data <= 8'hFF;
            15'd9819: data <= 8'hFF;
            15'd9820: data <= 8'hFF;
            15'd9821: data <= 8'hFF;
            15'd9822: data <= 8'hFC;
            15'd9823: data <= 8'hC0;
            15'd9824: data <= 8'h7F;
            15'd9825: data <= 8'hE0;
            15'd9826: data <= 8'h03;
            15'd9827: data <= 8'hFF;
            15'd9828: data <= 8'hF3;
            15'd9829: data <= 8'hFF;
            15'd9830: data <= 8'hFF;
            15'd9831: data <= 8'hFF;
            15'd9832: data <= 8'hFF;
            15'd9833: data <= 8'hFF;
            15'd9834: data <= 8'hFF;
            15'd9835: data <= 8'h80;
            15'd9836: data <= 8'h00;
            15'd9837: data <= 8'h00;
            15'd9838: data <= 8'h00;
            15'd9839: data <= 8'h00;
            15'd9840: data <= 8'h00;
            15'd9841: data <= 8'h00;
            15'd9842: data <= 8'h00;
            15'd9843: data <= 8'h00;
            15'd9844: data <= 8'h01;
            15'd9845: data <= 8'hFF;
            15'd9846: data <= 8'hFF;
            15'd9847: data <= 8'hFF;
            15'd9848: data <= 8'hFF;
            15'd9849: data <= 8'hFF;
            15'd9850: data <= 8'hFF;
            15'd9851: data <= 8'hFF;
            15'd9852: data <= 8'hF8;
            15'd9853: data <= 8'h00;
            15'd9854: data <= 8'h7F;
            15'd9855: data <= 8'hC7;
            15'd9856: data <= 8'hFF;
            15'd9857: data <= 8'hFF;
            15'd9858: data <= 8'hF1;
            15'd9859: data <= 8'hFF;
            15'd9860: data <= 8'hFF;
            15'd9861: data <= 8'hFF;
            15'd9862: data <= 8'hFF;
            15'd9863: data <= 8'hFF;
            15'd9864: data <= 8'hFF;
            15'd9865: data <= 8'h80;
            15'd9866: data <= 8'h00;
            15'd9867: data <= 8'h00;
            15'd9868: data <= 8'h00;
            15'd9869: data <= 8'h00;
            15'd9870: data <= 8'h00;
            15'd9871: data <= 8'h00;
            15'd9872: data <= 8'h00;
            15'd9873: data <= 8'h00;
            15'd9874: data <= 8'h01;
            15'd9875: data <= 8'hFF;
            15'd9876: data <= 8'hFF;
            15'd9877: data <= 8'hFF;
            15'd9878: data <= 8'hFF;
            15'd9879: data <= 8'hFF;
            15'd9880: data <= 8'hFF;
            15'd9881: data <= 8'hFF;
            15'd9882: data <= 8'hF8;
            15'd9883: data <= 8'h00;
            15'd9884: data <= 8'hFF;
            15'd9885: data <= 8'h80;
            15'd9886: data <= 8'h03;
            15'd9887: data <= 8'hFF;
            15'd9888: data <= 8'hE1;
            15'd9889: data <= 8'hFF;
            15'd9890: data <= 8'hFF;
            15'd9891: data <= 8'hFF;
            15'd9892: data <= 8'hFF;
            15'd9893: data <= 8'hFF;
            15'd9894: data <= 8'hFF;
            15'd9895: data <= 8'h80;
            15'd9896: data <= 8'h00;
            15'd9897: data <= 8'h00;
            15'd9898: data <= 8'h00;
            15'd9899: data <= 8'h00;
            15'd9900: data <= 8'h00;
            15'd9901: data <= 8'h00;
            15'd9902: data <= 8'h00;
            15'd9903: data <= 8'h00;
            15'd9904: data <= 8'h01;
            15'd9905: data <= 8'hFF;
            15'd9906: data <= 8'hFF;
            15'd9907: data <= 8'hFF;
            15'd9908: data <= 8'hFF;
            15'd9909: data <= 8'hFF;
            15'd9910: data <= 8'hFF;
            15'd9911: data <= 8'hFF;
            15'd9912: data <= 8'hF8;
            15'd9913: data <= 8'hC7;
            15'd9914: data <= 8'hFF;
            15'd9915: data <= 8'h88;
            15'd9916: data <= 8'h03;
            15'd9917: data <= 8'hFF;
            15'd9918: data <= 8'hE3;
            15'd9919: data <= 8'hFF;
            15'd9920: data <= 8'hFF;
            15'd9921: data <= 8'hFF;
            15'd9922: data <= 8'hFF;
            15'd9923: data <= 8'hFF;
            15'd9924: data <= 8'hFF;
            15'd9925: data <= 8'h80;
            15'd9926: data <= 8'h00;
            15'd9927: data <= 8'h00;
            15'd9928: data <= 8'h00;
            15'd9929: data <= 8'h00;
            15'd9930: data <= 8'h00;
            15'd9931: data <= 8'h00;
            15'd9932: data <= 8'h00;
            15'd9933: data <= 8'h00;
            15'd9934: data <= 8'h01;
            15'd9935: data <= 8'hFF;
            15'd9936: data <= 8'hFF;
            15'd9937: data <= 8'hFF;
            15'd9938: data <= 8'hFF;
            15'd9939: data <= 8'hFF;
            15'd9940: data <= 8'hFF;
            15'd9941: data <= 8'hFF;
            15'd9942: data <= 8'hF1;
            15'd9943: data <= 8'h87;
            15'd9944: data <= 8'hFF;
            15'd9945: data <= 8'h9F;
            15'd9946: data <= 8'hFF;
            15'd9947: data <= 8'hFF;
            15'd9948: data <= 8'hE3;
            15'd9949: data <= 8'hFF;
            15'd9950: data <= 8'hFF;
            15'd9951: data <= 8'hFF;
            15'd9952: data <= 8'hFF;
            15'd9953: data <= 8'hFF;
            15'd9954: data <= 8'hFF;
            15'd9955: data <= 8'h80;
            15'd9956: data <= 8'h00;
            15'd9957: data <= 8'h00;
            15'd9958: data <= 8'h00;
            15'd9959: data <= 8'h00;
            15'd9960: data <= 8'h00;
            15'd9961: data <= 8'h00;
            15'd9962: data <= 8'h00;
            15'd9963: data <= 8'h00;
            15'd9964: data <= 8'h01;
            15'd9965: data <= 8'hFF;
            15'd9966: data <= 8'hFF;
            15'd9967: data <= 8'hFF;
            15'd9968: data <= 8'hFF;
            15'd9969: data <= 8'hFF;
            15'd9970: data <= 8'hFF;
            15'd9971: data <= 8'hFF;
            15'd9972: data <= 8'hF1;
            15'd9973: data <= 8'hC7;
            15'd9974: data <= 8'hFF;
            15'd9975: data <= 8'hF8;
            15'd9976: data <= 8'h01;
            15'd9977: data <= 8'hFF;
            15'd9978: data <= 8'hE3;
            15'd9979: data <= 8'hFF;
            15'd9980: data <= 8'hFF;
            15'd9981: data <= 8'hFF;
            15'd9982: data <= 8'hFF;
            15'd9983: data <= 8'hFF;
            15'd9984: data <= 8'hFF;
            15'd9985: data <= 8'h80;
            15'd9986: data <= 8'h00;
            15'd9987: data <= 8'h00;
            15'd9988: data <= 8'h00;
            15'd9989: data <= 8'h00;
            15'd9990: data <= 8'h00;
            15'd9991: data <= 8'h00;
            15'd9992: data <= 8'h00;
            15'd9993: data <= 8'h00;
            15'd9994: data <= 8'h01;
            15'd9995: data <= 8'hFF;
            15'd9996: data <= 8'hFF;
            15'd9997: data <= 8'hFF;
            15'd9998: data <= 8'hFF;
            15'd9999: data <= 8'hFF;
            15'd10000: data <= 8'hFF;
            15'd10001: data <= 8'hFF;
            15'd10002: data <= 8'hF3;
            15'd10003: data <= 8'hC1;
            15'd10004: data <= 8'hFF;
            15'd10005: data <= 8'hF0;
            15'd10006: data <= 8'h01;
            15'd10007: data <= 8'hFF;
            15'd10008: data <= 8'hF3;
            15'd10009: data <= 8'hFF;
            15'd10010: data <= 8'hFF;
            15'd10011: data <= 8'hFF;
            15'd10012: data <= 8'hFF;
            15'd10013: data <= 8'hFF;
            15'd10014: data <= 8'hFF;
            15'd10015: data <= 8'h80;
            15'd10016: data <= 8'h00;
            15'd10017: data <= 8'h00;
            15'd10018: data <= 8'h00;
            15'd10019: data <= 8'h00;
            15'd10020: data <= 8'h00;
            15'd10021: data <= 8'h00;
            15'd10022: data <= 8'h00;
            15'd10023: data <= 8'h00;
            15'd10024: data <= 8'h01;
            15'd10025: data <= 8'hFF;
            15'd10026: data <= 8'hFF;
            15'd10027: data <= 8'hFF;
            15'd10028: data <= 8'hFF;
            15'd10029: data <= 8'hFF;
            15'd10030: data <= 8'hFF;
            15'd10031: data <= 8'hFF;
            15'd10032: data <= 8'hFE;
            15'd10033: data <= 8'h00;
            15'd10034: data <= 8'h7F;
            15'd10035: data <= 8'hF8;
            15'd10036: data <= 8'h11;
            15'd10037: data <= 8'hFF;
            15'd10038: data <= 8'hF3;
            15'd10039: data <= 8'hFF;
            15'd10040: data <= 8'hFF;
            15'd10041: data <= 8'hFF;
            15'd10042: data <= 8'hFF;
            15'd10043: data <= 8'hFF;
            15'd10044: data <= 8'hFF;
            15'd10045: data <= 8'h80;
            15'd10046: data <= 8'h00;
            15'd10047: data <= 8'h00;
            15'd10048: data <= 8'h00;
            15'd10049: data <= 8'h00;
            15'd10050: data <= 8'h00;
            15'd10051: data <= 8'h00;
            15'd10052: data <= 8'h00;
            15'd10053: data <= 8'h00;
            15'd10054: data <= 8'h01;
            15'd10055: data <= 8'hFF;
            15'd10056: data <= 8'hFF;
            15'd10057: data <= 8'hFF;
            15'd10058: data <= 8'hFF;
            15'd10059: data <= 8'hFF;
            15'd10060: data <= 8'hFF;
            15'd10061: data <= 8'hFF;
            15'd10062: data <= 8'hFC;
            15'd10063: data <= 8'h00;
            15'd10064: data <= 8'h7F;
            15'd10065: data <= 8'hFF;
            15'd10066: data <= 8'hF9;
            15'd10067: data <= 8'hFF;
            15'd10068: data <= 8'hF3;
            15'd10069: data <= 8'hFF;
            15'd10070: data <= 8'hFF;
            15'd10071: data <= 8'hFF;
            15'd10072: data <= 8'hFF;
            15'd10073: data <= 8'hFF;
            15'd10074: data <= 8'hFF;
            15'd10075: data <= 8'h80;
            15'd10076: data <= 8'h00;
            15'd10077: data <= 8'h00;
            15'd10078: data <= 8'h00;
            15'd10079: data <= 8'h00;
            15'd10080: data <= 8'h00;
            15'd10081: data <= 8'h00;
            15'd10082: data <= 8'h00;
            15'd10083: data <= 8'h00;
            15'd10084: data <= 8'h01;
            15'd10085: data <= 8'hFF;
            15'd10086: data <= 8'hFF;
            15'd10087: data <= 8'hFF;
            15'd10088: data <= 8'hFF;
            15'd10089: data <= 8'hFF;
            15'd10090: data <= 8'hFF;
            15'd10091: data <= 8'hFF;
            15'd10092: data <= 8'hFE;
            15'd10093: data <= 8'h03;
            15'd10094: data <= 8'hFF;
            15'd10095: data <= 8'hFF;
            15'd10096: data <= 8'hF9;
            15'd10097: data <= 8'hFF;
            15'd10098: data <= 8'hFF;
            15'd10099: data <= 8'hFF;
            15'd10100: data <= 8'hFF;
            15'd10101: data <= 8'hFF;
            15'd10102: data <= 8'hFF;
            15'd10103: data <= 8'hFF;
            15'd10104: data <= 8'hFF;
            15'd10105: data <= 8'h80;
            15'd10106: data <= 8'h00;
            15'd10107: data <= 8'h00;
            15'd10108: data <= 8'h00;
            15'd10109: data <= 8'h00;
            15'd10110: data <= 8'h00;
            15'd10111: data <= 8'h00;
            15'd10112: data <= 8'h00;
            15'd10113: data <= 8'h00;
            15'd10114: data <= 8'h01;
            15'd10115: data <= 8'hFF;
            15'd10116: data <= 8'hFF;
            15'd10117: data <= 8'hFF;
            15'd10118: data <= 8'hFF;
            15'd10119: data <= 8'hFF;
            15'd10120: data <= 8'hFF;
            15'd10121: data <= 8'hFF;
            15'd10122: data <= 8'hFF;
            15'd10123: data <= 8'hC7;
            15'd10124: data <= 8'hFF;
            15'd10125: data <= 8'hFF;
            15'd10126: data <= 8'hF8;
            15'd10127: data <= 8'hFF;
            15'd10128: data <= 8'hFF;
            15'd10129: data <= 8'hFF;
            15'd10130: data <= 8'hFF;
            15'd10131: data <= 8'hFF;
            15'd10132: data <= 8'hFF;
            15'd10133: data <= 8'hFF;
            15'd10134: data <= 8'hFF;
            15'd10135: data <= 8'h80;
            15'd10136: data <= 8'h00;
            15'd10137: data <= 8'h00;
            15'd10138: data <= 8'h00;
            15'd10139: data <= 8'h00;
            15'd10140: data <= 8'h00;
            15'd10141: data <= 8'h00;
            15'd10142: data <= 8'h00;
            15'd10143: data <= 8'h00;
            15'd10144: data <= 8'h01;
            15'd10145: data <= 8'hFF;
            15'd10146: data <= 8'hFF;
            15'd10147: data <= 8'hFF;
            15'd10148: data <= 8'hFF;
            15'd10149: data <= 8'hFF;
            15'd10150: data <= 8'hFF;
            15'd10151: data <= 8'hFF;
            15'd10152: data <= 8'hFF;
            15'd10153: data <= 8'hC7;
            15'd10154: data <= 8'hFF;
            15'd10155: data <= 8'hFF;
            15'd10156: data <= 8'hF8;
            15'd10157: data <= 8'hBF;
            15'd10158: data <= 8'hE7;
            15'd10159: data <= 8'hFF;
            15'd10160: data <= 8'hFF;
            15'd10161: data <= 8'hFF;
            15'd10162: data <= 8'hFF;
            15'd10163: data <= 8'hFF;
            15'd10164: data <= 8'hFF;
            15'd10165: data <= 8'h80;
            15'd10166: data <= 8'h00;
            15'd10167: data <= 8'h00;
            15'd10168: data <= 8'h00;
            15'd10169: data <= 8'h00;
            15'd10170: data <= 8'h00;
            15'd10171: data <= 8'h00;
            15'd10172: data <= 8'h00;
            15'd10173: data <= 8'h00;
            15'd10174: data <= 8'h01;
            15'd10175: data <= 8'hFF;
            15'd10176: data <= 8'hFF;
            15'd10177: data <= 8'hFF;
            15'd10178: data <= 8'hFF;
            15'd10179: data <= 8'hFF;
            15'd10180: data <= 8'hFF;
            15'd10181: data <= 8'hFF;
            15'd10182: data <= 8'hF1;
            15'd10183: data <= 8'h00;
            15'd10184: data <= 8'h1F;
            15'd10185: data <= 8'hFF;
            15'd10186: data <= 8'hFC;
            15'd10187: data <= 8'h1F;
            15'd10188: data <= 8'hE3;
            15'd10189: data <= 8'hFF;
            15'd10190: data <= 8'hFF;
            15'd10191: data <= 8'hFF;
            15'd10192: data <= 8'hFF;
            15'd10193: data <= 8'hFF;
            15'd10194: data <= 8'hFF;
            15'd10195: data <= 8'h80;
            15'd10196: data <= 8'h00;
            15'd10197: data <= 8'h00;
            15'd10198: data <= 8'h00;
            15'd10199: data <= 8'h00;
            15'd10200: data <= 8'h00;
            15'd10201: data <= 8'h00;
            15'd10202: data <= 8'h00;
            15'd10203: data <= 8'h00;
            15'd10204: data <= 8'h01;
            15'd10205: data <= 8'hFF;
            15'd10206: data <= 8'hFF;
            15'd10207: data <= 8'hFF;
            15'd10208: data <= 8'hFF;
            15'd10209: data <= 8'hFF;
            15'd10210: data <= 8'hFF;
            15'd10211: data <= 8'hFF;
            15'd10212: data <= 8'hE0;
            15'd10213: data <= 8'h00;
            15'd10214: data <= 8'h0F;
            15'd10215: data <= 8'hFF;
            15'd10216: data <= 8'hFC;
            15'd10217: data <= 8'h1F;
            15'd10218: data <= 8'hE7;
            15'd10219: data <= 8'hFF;
            15'd10220: data <= 8'hFF;
            15'd10221: data <= 8'hFF;
            15'd10222: data <= 8'hFF;
            15'd10223: data <= 8'hFF;
            15'd10224: data <= 8'hFF;
            15'd10225: data <= 8'h80;
            15'd10226: data <= 8'h00;
            15'd10227: data <= 8'h00;
            15'd10228: data <= 8'h00;
            15'd10229: data <= 8'h00;
            15'd10230: data <= 8'h00;
            15'd10231: data <= 8'h00;
            15'd10232: data <= 8'h00;
            15'd10233: data <= 8'h00;
            15'd10234: data <= 8'h01;
            15'd10235: data <= 8'hFF;
            15'd10236: data <= 8'hFF;
            15'd10237: data <= 8'hFF;
            15'd10238: data <= 8'hFF;
            15'd10239: data <= 8'hFF;
            15'd10240: data <= 8'hFF;
            15'd10241: data <= 8'hFF;
            15'd10242: data <= 8'hE0;
            15'd10243: data <= 8'h00;
            15'd10244: data <= 8'h0F;
            15'd10245: data <= 8'hFF;
            15'd10246: data <= 8'hFE;
            15'd10247: data <= 8'h3F;
            15'd10248: data <= 8'hFF;
            15'd10249: data <= 8'hFF;
            15'd10250: data <= 8'hFF;
            15'd10251: data <= 8'hFF;
            15'd10252: data <= 8'hFF;
            15'd10253: data <= 8'hFF;
            15'd10254: data <= 8'hFF;
            15'd10255: data <= 8'h80;
            15'd10256: data <= 8'h00;
            15'd10257: data <= 8'h00;
            15'd10258: data <= 8'h00;
            15'd10259: data <= 8'h00;
            15'd10260: data <= 8'h00;
            15'd10261: data <= 8'h00;
            15'd10262: data <= 8'h00;
            15'd10263: data <= 8'h00;
            15'd10264: data <= 8'h01;
            15'd10265: data <= 8'hFF;
            15'd10266: data <= 8'hFF;
            15'd10267: data <= 8'hFF;
            15'd10268: data <= 8'hFF;
            15'd10269: data <= 8'hFF;
            15'd10270: data <= 8'hFF;
            15'd10271: data <= 8'hFF;
            15'd10272: data <= 8'hF7;
            15'd10273: data <= 8'hFF;
            15'd10274: data <= 8'hFF;
            15'd10275: data <= 8'hFF;
            15'd10276: data <= 8'hFF;
            15'd10277: data <= 8'hFF;
            15'd10278: data <= 8'hFF;
            15'd10279: data <= 8'hFF;
            15'd10280: data <= 8'hFF;
            15'd10281: data <= 8'hFF;
            15'd10282: data <= 8'hFF;
            15'd10283: data <= 8'hFF;
            15'd10284: data <= 8'hFF;
            15'd10285: data <= 8'h80;
            15'd10286: data <= 8'h00;
            15'd10287: data <= 8'h00;
            15'd10288: data <= 8'h00;
            15'd10289: data <= 8'h00;
            15'd10290: data <= 8'h00;
            15'd10291: data <= 8'h00;
            15'd10292: data <= 8'h00;
            15'd10293: data <= 8'h00;
            15'd10294: data <= 8'h01;
            15'd10295: data <= 8'hFF;
            15'd10296: data <= 8'hFF;
            15'd10297: data <= 8'hFF;
            15'd10298: data <= 8'hFF;
            15'd10299: data <= 8'hFF;
            15'd10300: data <= 8'hFF;
            15'd10301: data <= 8'hFF;
            15'd10302: data <= 8'hFF;
            15'd10303: data <= 8'hFF;
            15'd10304: data <= 8'hFF;
            15'd10305: data <= 8'hFF;
            15'd10306: data <= 8'hFF;
            15'd10307: data <= 8'hFF;
            15'd10308: data <= 8'hFF;
            15'd10309: data <= 8'hFF;
            15'd10310: data <= 8'hFF;
            15'd10311: data <= 8'hFF;
            15'd10312: data <= 8'hFF;
            15'd10313: data <= 8'hFF;
            15'd10314: data <= 8'hFF;
            15'd10315: data <= 8'h80;
            15'd10316: data <= 8'h00;
            15'd10317: data <= 8'h00;
            15'd10318: data <= 8'h00;
            15'd10319: data <= 8'h00;
            15'd10320: data <= 8'h00;
            15'd10321: data <= 8'h00;
            15'd10322: data <= 8'h00;
            15'd10323: data <= 8'h00;
            15'd10324: data <= 8'h01;
            15'd10325: data <= 8'hFF;
            15'd10326: data <= 8'hFF;
            15'd10327: data <= 8'hFF;
            15'd10328: data <= 8'hFF;
            15'd10329: data <= 8'hFF;
            15'd10330: data <= 8'hFF;
            15'd10331: data <= 8'hFF;
            15'd10332: data <= 8'hFF;
            15'd10333: data <= 8'hFF;
            15'd10334: data <= 8'hFF;
            15'd10335: data <= 8'hFF;
            15'd10336: data <= 8'hFF;
            15'd10337: data <= 8'hFF;
            15'd10338: data <= 8'hFF;
            15'd10339: data <= 8'hFF;
            15'd10340: data <= 8'hFF;
            15'd10341: data <= 8'hFF;
            15'd10342: data <= 8'hFF;
            15'd10343: data <= 8'hFF;
            15'd10344: data <= 8'hFF;
            15'd10345: data <= 8'h80;
            15'd10346: data <= 8'h00;
            15'd10347: data <= 8'h00;
            15'd10348: data <= 8'h00;
            15'd10349: data <= 8'h00;
            15'd10350: data <= 8'h00;
            15'd10351: data <= 8'h00;
            15'd10352: data <= 8'h00;
            15'd10353: data <= 8'h00;
            15'd10354: data <= 8'h01;
            15'd10355: data <= 8'hFF;
            15'd10356: data <= 8'hFF;
            15'd10357: data <= 8'hFF;
            15'd10358: data <= 8'hFF;
            15'd10359: data <= 8'hFF;
            15'd10360: data <= 8'hFF;
            15'd10361: data <= 8'hFF;
            15'd10362: data <= 8'hFF;
            15'd10363: data <= 8'hFF;
            15'd10364: data <= 8'hFF;
            15'd10365: data <= 8'hFF;
            15'd10366: data <= 8'hFF;
            15'd10367: data <= 8'hFF;
            15'd10368: data <= 8'hFF;
            15'd10369: data <= 8'hFF;
            15'd10370: data <= 8'hFF;
            15'd10371: data <= 8'hFF;
            15'd10372: data <= 8'hFF;
            15'd10373: data <= 8'hFF;
            15'd10374: data <= 8'hFF;
            15'd10375: data <= 8'h80;
            15'd10376: data <= 8'h00;
            15'd10377: data <= 8'h00;
            15'd10378: data <= 8'h00;
            15'd10379: data <= 8'h00;
            15'd10380: data <= 8'h00;
            15'd10381: data <= 8'h00;
            15'd10382: data <= 8'h00;
            15'd10383: data <= 8'h00;
            15'd10384: data <= 8'h01;
            15'd10385: data <= 8'hFF;
            15'd10386: data <= 8'hFF;
            15'd10387: data <= 8'hFF;
            15'd10388: data <= 8'hFF;
            15'd10389: data <= 8'hFF;
            15'd10390: data <= 8'hFF;
            15'd10391: data <= 8'hFF;
            15'd10392: data <= 8'hFF;
            15'd10393: data <= 8'hFF;
            15'd10394: data <= 8'hFF;
            15'd10395: data <= 8'hFF;
            15'd10396: data <= 8'hFF;
            15'd10397: data <= 8'hFF;
            15'd10398: data <= 8'hFF;
            15'd10399: data <= 8'hFF;
            15'd10400: data <= 8'hFF;
            15'd10401: data <= 8'hFF;
            15'd10402: data <= 8'hFF;
            15'd10403: data <= 8'hFF;
            15'd10404: data <= 8'hFF;
            15'd10405: data <= 8'h80;
            15'd10406: data <= 8'h00;
            15'd10407: data <= 8'h00;
            15'd10408: data <= 8'h00;
            15'd10409: data <= 8'h00;
            15'd10410: data <= 8'h00;
            15'd10411: data <= 8'h00;
            15'd10412: data <= 8'h00;
            15'd10413: data <= 8'h00;
            15'd10414: data <= 8'h01;
            15'd10415: data <= 8'hFF;
            15'd10416: data <= 8'hFF;
            15'd10417: data <= 8'hFF;
            15'd10418: data <= 8'hFF;
            15'd10419: data <= 8'hFF;
            15'd10420: data <= 8'hFF;
            15'd10421: data <= 8'hFF;
            15'd10422: data <= 8'hFF;
            15'd10423: data <= 8'hFF;
            15'd10424: data <= 8'hFF;
            15'd10425: data <= 8'hFF;
            15'd10426: data <= 8'hFF;
            15'd10427: data <= 8'hFF;
            15'd10428: data <= 8'hFF;
            15'd10429: data <= 8'hFF;
            15'd10430: data <= 8'hFF;
            15'd10431: data <= 8'hFF;
            15'd10432: data <= 8'hFF;
            15'd10433: data <= 8'hFF;
            15'd10434: data <= 8'hFF;
            15'd10435: data <= 8'h80;
            15'd10436: data <= 8'h00;
            15'd10437: data <= 8'h00;
            15'd10438: data <= 8'h00;
            15'd10439: data <= 8'h00;
            15'd10440: data <= 8'h00;
            15'd10441: data <= 8'h00;
            15'd10442: data <= 8'h00;
            15'd10443: data <= 8'h00;
            15'd10444: data <= 8'h01;
            15'd10445: data <= 8'hFF;
            15'd10446: data <= 8'hFF;
            15'd10447: data <= 8'hFF;
            15'd10448: data <= 8'hFF;
            15'd10449: data <= 8'hFF;
            15'd10450: data <= 8'hFF;
            15'd10451: data <= 8'hFF;
            15'd10452: data <= 8'hFF;
            15'd10453: data <= 8'hFF;
            15'd10454: data <= 8'hFF;
            15'd10455: data <= 8'hFF;
            15'd10456: data <= 8'hFF;
            15'd10457: data <= 8'hFF;
            15'd10458: data <= 8'hFF;
            15'd10459: data <= 8'hFF;
            15'd10460: data <= 8'hFF;
            15'd10461: data <= 8'hFF;
            15'd10462: data <= 8'hFF;
            15'd10463: data <= 8'hFF;
            15'd10464: data <= 8'hFF;
            15'd10465: data <= 8'h80;
            15'd10466: data <= 8'h00;
            15'd10467: data <= 8'h00;
            15'd10468: data <= 8'h00;
            15'd10469: data <= 8'h00;
            15'd10470: data <= 8'h00;
            15'd10471: data <= 8'h00;
            15'd10472: data <= 8'h00;
            15'd10473: data <= 8'h00;
            15'd10474: data <= 8'h01;
            15'd10475: data <= 8'hFF;
            15'd10476: data <= 8'hFF;
            15'd10477: data <= 8'hFF;
            15'd10478: data <= 8'hFF;
            15'd10479: data <= 8'hFF;
            15'd10480: data <= 8'hFF;
            15'd10481: data <= 8'hFF;
            15'd10482: data <= 8'hFF;
            15'd10483: data <= 8'hFF;
            15'd10484: data <= 8'hFF;
            15'd10485: data <= 8'hFF;
            15'd10486: data <= 8'hFF;
            15'd10487: data <= 8'hFF;
            15'd10488: data <= 8'hFF;
            15'd10489: data <= 8'hFF;
            15'd10490: data <= 8'hFF;
            15'd10491: data <= 8'hFF;
            15'd10492: data <= 8'hFF;
            15'd10493: data <= 8'hFF;
            15'd10494: data <= 8'hFF;
            15'd10495: data <= 8'h80;
            15'd10496: data <= 8'h00;
            15'd10497: data <= 8'h00;
            15'd10498: data <= 8'h00;
            15'd10499: data <= 8'h00;
            15'd10500: data <= 8'h00;
            15'd10501: data <= 8'h00;
            15'd10502: data <= 8'h00;
            15'd10503: data <= 8'h00;
            15'd10504: data <= 8'h01;
            15'd10505: data <= 8'hFF;
            15'd10506: data <= 8'hFF;
            15'd10507: data <= 8'hFF;
            15'd10508: data <= 8'hFF;
            15'd10509: data <= 8'hFF;
            15'd10510: data <= 8'hFF;
            15'd10511: data <= 8'hFF;
            15'd10512: data <= 8'hFF;
            15'd10513: data <= 8'hFF;
            15'd10514: data <= 8'hFF;
            15'd10515: data <= 8'hFF;
            15'd10516: data <= 8'hFF;
            15'd10517: data <= 8'hFF;
            15'd10518: data <= 8'hFF;
            15'd10519: data <= 8'hFF;
            15'd10520: data <= 8'hFF;
            15'd10521: data <= 8'hFF;
            15'd10522: data <= 8'hFF;
            15'd10523: data <= 8'hFF;
            15'd10524: data <= 8'hFF;
            15'd10525: data <= 8'h80;
            15'd10526: data <= 8'h00;
            15'd10527: data <= 8'h00;
            15'd10528: data <= 8'h00;
            15'd10529: data <= 8'h00;
            15'd10530: data <= 8'h00;
            15'd10531: data <= 8'h00;
            15'd10532: data <= 8'h00;
            15'd10533: data <= 8'h00;
            15'd10534: data <= 8'h01;
            15'd10535: data <= 8'hFF;
            15'd10536: data <= 8'hFF;
            15'd10537: data <= 8'hFF;
            15'd10538: data <= 8'hFF;
            15'd10539: data <= 8'hFF;
            15'd10540: data <= 8'hFF;
            15'd10541: data <= 8'hFF;
            15'd10542: data <= 8'hFF;
            15'd10543: data <= 8'hFF;
            15'd10544: data <= 8'hFF;
            15'd10545: data <= 8'hFF;
            15'd10546: data <= 8'hFF;
            15'd10547: data <= 8'hFF;
            15'd10548: data <= 8'hFF;
            15'd10549: data <= 8'hFF;
            15'd10550: data <= 8'hFF;
            15'd10551: data <= 8'hFF;
            15'd10552: data <= 8'hFF;
            15'd10553: data <= 8'hFF;
            15'd10554: data <= 8'hFF;
            15'd10555: data <= 8'h80;
            15'd10556: data <= 8'h00;
            15'd10557: data <= 8'h00;
            15'd10558: data <= 8'h00;
            15'd10559: data <= 8'h00;
            15'd10560: data <= 8'h00;
            15'd10561: data <= 8'h00;
            15'd10562: data <= 8'h00;
            15'd10563: data <= 8'h00;
            15'd10564: data <= 8'h01;
            15'd10565: data <= 8'hFF;
            15'd10566: data <= 8'hFF;
            15'd10567: data <= 8'hFF;
            15'd10568: data <= 8'hFF;
            15'd10569: data <= 8'hFF;
            15'd10570: data <= 8'hFF;
            15'd10571: data <= 8'hFF;
            15'd10572: data <= 8'hFF;
            15'd10573: data <= 8'hFF;
            15'd10574: data <= 8'hFF;
            15'd10575: data <= 8'hFF;
            15'd10576: data <= 8'hFF;
            15'd10577: data <= 8'hFF;
            15'd10578: data <= 8'hFF;
            15'd10579: data <= 8'hFF;
            15'd10580: data <= 8'hFF;
            15'd10581: data <= 8'hFF;
            15'd10582: data <= 8'hFF;
            15'd10583: data <= 8'hFF;
            15'd10584: data <= 8'hFF;
            15'd10585: data <= 8'h80;
            15'd10586: data <= 8'h00;
            15'd10587: data <= 8'h00;
            15'd10588: data <= 8'h00;
            15'd10589: data <= 8'h00;
            15'd10590: data <= 8'h00;
            15'd10591: data <= 8'h00;
            15'd10592: data <= 8'h00;
            15'd10593: data <= 8'h00;
            15'd10594: data <= 8'h01;
            15'd10595: data <= 8'hFF;
            15'd10596: data <= 8'hFF;
            15'd10597: data <= 8'hFF;
            15'd10598: data <= 8'hFF;
            15'd10599: data <= 8'hFF;
            15'd10600: data <= 8'hFF;
            15'd10601: data <= 8'hFF;
            15'd10602: data <= 8'hFF;
            15'd10603: data <= 8'hFF;
            15'd10604: data <= 8'hFF;
            15'd10605: data <= 8'hFF;
            15'd10606: data <= 8'hFF;
            15'd10607: data <= 8'hFF;
            15'd10608: data <= 8'hFF;
            15'd10609: data <= 8'hFF;
            15'd10610: data <= 8'hFF;
            15'd10611: data <= 8'hFF;
            15'd10612: data <= 8'hFF;
            15'd10613: data <= 8'hFF;
            15'd10614: data <= 8'hFF;
            15'd10615: data <= 8'h80;
            15'd10616: data <= 8'h00;
            15'd10617: data <= 8'h00;
            15'd10618: data <= 8'h00;
            15'd10619: data <= 8'h00;
            15'd10620: data <= 8'h00;
            15'd10621: data <= 8'h00;
            15'd10622: data <= 8'h00;
            15'd10623: data <= 8'h00;
            15'd10624: data <= 8'h01;
            15'd10625: data <= 8'hFF;
            15'd10626: data <= 8'hFF;
            15'd10627: data <= 8'hFF;
            15'd10628: data <= 8'hFF;
            15'd10629: data <= 8'hFF;
            15'd10630: data <= 8'hFF;
            15'd10631: data <= 8'hFF;
            15'd10632: data <= 8'hFF;
            15'd10633: data <= 8'hFF;
            15'd10634: data <= 8'hFF;
            15'd10635: data <= 8'hFF;
            15'd10636: data <= 8'hFF;
            15'd10637: data <= 8'hFF;
            15'd10638: data <= 8'hFF;
            15'd10639: data <= 8'hFF;
            15'd10640: data <= 8'hFF;
            15'd10641: data <= 8'hFF;
            15'd10642: data <= 8'hFF;
            15'd10643: data <= 8'hFF;
            15'd10644: data <= 8'hFF;
            15'd10645: data <= 8'h80;
            15'd10646: data <= 8'h00;
            15'd10647: data <= 8'h00;
            15'd10648: data <= 8'h00;
            15'd10649: data <= 8'h00;
            15'd10650: data <= 8'h00;
            15'd10651: data <= 8'h00;
            15'd10652: data <= 8'h00;
            15'd10653: data <= 8'h00;
            15'd10654: data <= 8'h01;
            15'd10655: data <= 8'hFF;
            15'd10656: data <= 8'hFF;
            15'd10657: data <= 8'hFF;
            15'd10658: data <= 8'hFF;
            15'd10659: data <= 8'hFF;
            15'd10660: data <= 8'hFF;
            15'd10661: data <= 8'hFF;
            15'd10662: data <= 8'hFF;
            15'd10663: data <= 8'hFF;
            15'd10664: data <= 8'hFF;
            15'd10665: data <= 8'hFF;
            15'd10666: data <= 8'hFF;
            15'd10667: data <= 8'hFF;
            15'd10668: data <= 8'hFF;
            15'd10669: data <= 8'hFF;
            15'd10670: data <= 8'hFF;
            15'd10671: data <= 8'hFF;
            15'd10672: data <= 8'hFF;
            15'd10673: data <= 8'hFF;
            15'd10674: data <= 8'hFF;
            15'd10675: data <= 8'h80;
            15'd10676: data <= 8'h00;
            15'd10677: data <= 8'h00;
            15'd10678: data <= 8'h00;
            15'd10679: data <= 8'h00;
            15'd10680: data <= 8'h00;
            15'd10681: data <= 8'h00;
            15'd10682: data <= 8'h00;
            15'd10683: data <= 8'h00;
            15'd10684: data <= 8'h01;
            15'd10685: data <= 8'hFF;
            15'd10686: data <= 8'hFF;
            15'd10687: data <= 8'hFF;
            15'd10688: data <= 8'hFF;
            15'd10689: data <= 8'hFF;
            15'd10690: data <= 8'hFF;
            15'd10691: data <= 8'hFF;
            15'd10692: data <= 8'hFF;
            15'd10693: data <= 8'hFF;
            15'd10694: data <= 8'hFF;
            15'd10695: data <= 8'hFF;
            15'd10696: data <= 8'hFF;
            15'd10697: data <= 8'hFF;
            15'd10698: data <= 8'hFF;
            15'd10699: data <= 8'hFF;
            15'd10700: data <= 8'hFF;
            15'd10701: data <= 8'hFF;
            15'd10702: data <= 8'hFF;
            15'd10703: data <= 8'hFF;
            15'd10704: data <= 8'hFF;
            15'd10705: data <= 8'h80;
            15'd10706: data <= 8'h00;
            15'd10707: data <= 8'h00;
            15'd10708: data <= 8'h00;
            15'd10709: data <= 8'h00;
            15'd10710: data <= 8'h00;
            15'd10711: data <= 8'h00;
            15'd10712: data <= 8'h00;
            15'd10713: data <= 8'h00;
            15'd10714: data <= 8'h01;
            15'd10715: data <= 8'hFF;
            15'd10716: data <= 8'hFF;
            15'd10717: data <= 8'hFF;
            15'd10718: data <= 8'hFF;
            15'd10719: data <= 8'hFF;
            15'd10720: data <= 8'hFF;
            15'd10721: data <= 8'hFF;
            15'd10722: data <= 8'hFF;
            15'd10723: data <= 8'hFF;
            15'd10724: data <= 8'hFF;
            15'd10725: data <= 8'hFF;
            15'd10726: data <= 8'hFF;
            15'd10727: data <= 8'hFF;
            15'd10728: data <= 8'hFF;
            15'd10729: data <= 8'hFF;
            15'd10730: data <= 8'hFF;
            15'd10731: data <= 8'hFF;
            15'd10732: data <= 8'hFF;
            15'd10733: data <= 8'hFF;
            15'd10734: data <= 8'hFF;
            15'd10735: data <= 8'h80;
            15'd10736: data <= 8'h00;
            15'd10737: data <= 8'h00;
            15'd10738: data <= 8'h00;
            15'd10739: data <= 8'h00;
            15'd10740: data <= 8'h00;
            15'd10741: data <= 8'h00;
            15'd10742: data <= 8'h00;
            15'd10743: data <= 8'h00;
            15'd10744: data <= 8'h01;
            15'd10745: data <= 8'hFF;
            15'd10746: data <= 8'hFF;
            15'd10747: data <= 8'hFF;
            15'd10748: data <= 8'hFF;
            15'd10749: data <= 8'hFF;
            15'd10750: data <= 8'hFF;
            15'd10751: data <= 8'hFF;
            15'd10752: data <= 8'hFF;
            15'd10753: data <= 8'hFF;
            15'd10754: data <= 8'hFF;
            15'd10755: data <= 8'hFF;
            15'd10756: data <= 8'hFF;
            15'd10757: data <= 8'hFF;
            15'd10758: data <= 8'hFF;
            15'd10759: data <= 8'hFF;
            15'd10760: data <= 8'hFF;
            15'd10761: data <= 8'hFF;
            15'd10762: data <= 8'hFF;
            15'd10763: data <= 8'hFF;
            15'd10764: data <= 8'hFF;
            15'd10765: data <= 8'h80;
            15'd10766: data <= 8'h00;
            15'd10767: data <= 8'h00;
            15'd10768: data <= 8'h00;
            15'd10769: data <= 8'h00;
            15'd10770: data <= 8'h00;
            15'd10771: data <= 8'h00;
            15'd10772: data <= 8'h00;
            15'd10773: data <= 8'h00;
            15'd10774: data <= 8'h01;
            15'd10775: data <= 8'hFF;
            15'd10776: data <= 8'hFF;
            15'd10777: data <= 8'hFF;
            15'd10778: data <= 8'hFF;
            15'd10779: data <= 8'hFF;
            15'd10780: data <= 8'hFF;
            15'd10781: data <= 8'hFF;
            15'd10782: data <= 8'hFF;
            15'd10783: data <= 8'hFF;
            15'd10784: data <= 8'hFF;
            15'd10785: data <= 8'hFF;
            15'd10786: data <= 8'hFF;
            15'd10787: data <= 8'hFF;
            15'd10788: data <= 8'hFF;
            15'd10789: data <= 8'hFF;
            15'd10790: data <= 8'hFF;
            15'd10791: data <= 8'hFF;
            15'd10792: data <= 8'hFF;
            15'd10793: data <= 8'hFF;
            15'd10794: data <= 8'hFF;
            15'd10795: data <= 8'h80;
            15'd10796: data <= 8'h00;
            15'd10797: data <= 8'h00;
            15'd10798: data <= 8'h00;
            15'd10799: data <= 8'h00;
            15'd10800: data <= 8'h00;
            15'd10801: data <= 8'h00;
            15'd10802: data <= 8'h00;
            15'd10803: data <= 8'h00;
            15'd10804: data <= 8'h00;
            15'd10805: data <= 8'h03;
            15'd10806: data <= 8'hFF;
            15'd10807: data <= 8'hFF;
            15'd10808: data <= 8'hFF;
            15'd10809: data <= 8'hFF;
            15'd10810: data <= 8'hFF;
            15'd10811: data <= 8'hFF;
            15'd10812: data <= 8'hFF;
            15'd10813: data <= 8'hFF;
            15'd10814: data <= 8'hFF;
            15'd10815: data <= 8'hFF;
            15'd10816: data <= 8'hFF;
            15'd10817: data <= 8'hFF;
            15'd10818: data <= 8'hFF;
            15'd10819: data <= 8'hFF;
            15'd10820: data <= 8'hFF;
            15'd10821: data <= 8'hFF;
            15'd10822: data <= 8'hFF;
            15'd10823: data <= 8'hFF;
            15'd10824: data <= 8'h80;
            15'd10825: data <= 8'h00;
            15'd10826: data <= 8'h00;
            15'd10827: data <= 8'h00;
            15'd10828: data <= 8'h00;
            15'd10829: data <= 8'h00;
            15'd10830: data <= 8'h00;
            15'd10831: data <= 8'h00;
            15'd10832: data <= 8'h00;
            15'd10833: data <= 8'h00;
            15'd10834: data <= 8'h00;
            15'd10835: data <= 8'h03;
            15'd10836: data <= 8'hFF;
            15'd10837: data <= 8'hFF;
            15'd10838: data <= 8'hFF;
            15'd10839: data <= 8'hFF;
            15'd10840: data <= 8'hFF;
            15'd10841: data <= 8'hFF;
            15'd10842: data <= 8'hFF;
            15'd10843: data <= 8'hFF;
            15'd10844: data <= 8'hFF;
            15'd10845: data <= 8'hFF;
            15'd10846: data <= 8'hFF;
            15'd10847: data <= 8'hFF;
            15'd10848: data <= 8'hFF;
            15'd10849: data <= 8'hFF;
            15'd10850: data <= 8'hFF;
            15'd10851: data <= 8'hFF;
            15'd10852: data <= 8'hFF;
            15'd10853: data <= 8'hFF;
            15'd10854: data <= 8'h80;
            15'd10855: data <= 8'h00;
            15'd10856: data <= 8'h00;
            15'd10857: data <= 8'h00;
            15'd10858: data <= 8'h00;
            15'd10859: data <= 8'h00;
            15'd10860: data <= 8'h00;
            15'd10861: data <= 8'h00;
            15'd10862: data <= 8'h00;
            15'd10863: data <= 8'h00;
            15'd10864: data <= 8'h00;
            15'd10865: data <= 8'h03;
            15'd10866: data <= 8'hFF;
            15'd10867: data <= 8'hFF;
            15'd10868: data <= 8'hFF;
            15'd10869: data <= 8'hFF;
            15'd10870: data <= 8'hFF;
            15'd10871: data <= 8'hFF;
            15'd10872: data <= 8'hFF;
            15'd10873: data <= 8'hFF;
            15'd10874: data <= 8'hFF;
            15'd10875: data <= 8'hFF;
            15'd10876: data <= 8'hFF;
            15'd10877: data <= 8'hFF;
            15'd10878: data <= 8'hFF;
            15'd10879: data <= 8'hFF;
            15'd10880: data <= 8'hFF;
            15'd10881: data <= 8'hFF;
            15'd10882: data <= 8'hFF;
            15'd10883: data <= 8'hFF;
            15'd10884: data <= 8'h80;
            15'd10885: data <= 8'h00;
            15'd10886: data <= 8'h00;
            15'd10887: data <= 8'h00;
            15'd10888: data <= 8'h00;
            15'd10889: data <= 8'h00;
            15'd10890: data <= 8'h00;
            15'd10891: data <= 8'h00;
            15'd10892: data <= 8'h00;
            15'd10893: data <= 8'h00;
            15'd10894: data <= 8'h00;
            15'd10895: data <= 8'h03;
            15'd10896: data <= 8'hFF;
            15'd10897: data <= 8'hFF;
            15'd10898: data <= 8'hFF;
            15'd10899: data <= 8'hFF;
            15'd10900: data <= 8'hFF;
            15'd10901: data <= 8'hFF;
            15'd10902: data <= 8'hFF;
            15'd10903: data <= 8'hFF;
            15'd10904: data <= 8'hFF;
            15'd10905: data <= 8'hFF;
            15'd10906: data <= 8'hFF;
            15'd10907: data <= 8'hFF;
            15'd10908: data <= 8'hFF;
            15'd10909: data <= 8'hFF;
            15'd10910: data <= 8'hFF;
            15'd10911: data <= 8'hFF;
            15'd10912: data <= 8'hFF;
            15'd10913: data <= 8'hFF;
            15'd10914: data <= 8'h80;
            15'd10915: data <= 8'h00;
            15'd10916: data <= 8'h00;
            15'd10917: data <= 8'h00;
            15'd10918: data <= 8'h00;
            15'd10919: data <= 8'h00;
            15'd10920: data <= 8'h00;
            15'd10921: data <= 8'h00;
            15'd10922: data <= 8'h00;
            15'd10923: data <= 8'h00;
            15'd10924: data <= 8'h00;
            15'd10925: data <= 8'h03;
            15'd10926: data <= 8'hFF;
            15'd10927: data <= 8'hFF;
            15'd10928: data <= 8'hFF;
            15'd10929: data <= 8'hFF;
            15'd10930: data <= 8'hFF;
            15'd10931: data <= 8'hFF;
            15'd10932: data <= 8'hFF;
            15'd10933: data <= 8'hFF;
            15'd10934: data <= 8'hFF;
            15'd10935: data <= 8'hFF;
            15'd10936: data <= 8'hFF;
            15'd10937: data <= 8'hFF;
            15'd10938: data <= 8'hFF;
            15'd10939: data <= 8'hFF;
            15'd10940: data <= 8'hFF;
            15'd10941: data <= 8'hFF;
            15'd10942: data <= 8'hFF;
            15'd10943: data <= 8'hFF;
            15'd10944: data <= 8'h80;
            15'd10945: data <= 8'h00;
            15'd10946: data <= 8'h00;
            15'd10947: data <= 8'h00;
            15'd10948: data <= 8'h00;
            15'd10949: data <= 8'h00;
            15'd10950: data <= 8'h00;
            15'd10951: data <= 8'h00;
            15'd10952: data <= 8'h00;
            15'd10953: data <= 8'h00;
            15'd10954: data <= 8'h00;
            15'd10955: data <= 8'h03;
            15'd10956: data <= 8'hFF;
            15'd10957: data <= 8'hFF;
            15'd10958: data <= 8'hFF;
            15'd10959: data <= 8'hFF;
            15'd10960: data <= 8'hFF;
            15'd10961: data <= 8'hFF;
            15'd10962: data <= 8'hFF;
            15'd10963: data <= 8'hFF;
            15'd10964: data <= 8'hFF;
            15'd10965: data <= 8'hFF;
            15'd10966: data <= 8'hFF;
            15'd10967: data <= 8'hFF;
            15'd10968: data <= 8'hFF;
            15'd10969: data <= 8'hFF;
            15'd10970: data <= 8'hFF;
            15'd10971: data <= 8'hFF;
            15'd10972: data <= 8'hFF;
            15'd10973: data <= 8'hFF;
            15'd10974: data <= 8'h80;
            15'd10975: data <= 8'h00;
            15'd10976: data <= 8'h00;
            15'd10977: data <= 8'h00;
            15'd10978: data <= 8'h00;
            15'd10979: data <= 8'h00;
            15'd10980: data <= 8'h00;
            15'd10981: data <= 8'h00;
            15'd10982: data <= 8'h00;
            15'd10983: data <= 8'h00;
            15'd10984: data <= 8'h00;
            15'd10985: data <= 8'h03;
            15'd10986: data <= 8'hFF;
            15'd10987: data <= 8'hFF;
            15'd10988: data <= 8'hFF;
            15'd10989: data <= 8'hFF;
            15'd10990: data <= 8'hFF;
            15'd10991: data <= 8'hFF;
            15'd10992: data <= 8'hFF;
            15'd10993: data <= 8'hFF;
            15'd10994: data <= 8'hFF;
            15'd10995: data <= 8'hFF;
            15'd10996: data <= 8'hFF;
            15'd10997: data <= 8'hFF;
            15'd10998: data <= 8'hFF;
            15'd10999: data <= 8'hFF;
            15'd11000: data <= 8'hFF;
            15'd11001: data <= 8'hFF;
            15'd11002: data <= 8'hFF;
            15'd11003: data <= 8'hFF;
            15'd11004: data <= 8'h80;
            15'd11005: data <= 8'h00;
            15'd11006: data <= 8'h00;
            15'd11007: data <= 8'h00;
            15'd11008: data <= 8'h00;
            15'd11009: data <= 8'h00;
            15'd11010: data <= 8'h00;
            15'd11011: data <= 8'h00;
            15'd11012: data <= 8'h00;
            15'd11013: data <= 8'h00;
            15'd11014: data <= 8'h00;
            15'd11015: data <= 8'h03;
            15'd11016: data <= 8'hFF;
            15'd11017: data <= 8'hFF;
            15'd11018: data <= 8'hFF;
            15'd11019: data <= 8'hFF;
            15'd11020: data <= 8'hFF;
            15'd11021: data <= 8'hFF;
            15'd11022: data <= 8'hFF;
            15'd11023: data <= 8'hFF;
            15'd11024: data <= 8'hFF;
            15'd11025: data <= 8'hFF;
            15'd11026: data <= 8'hFF;
            15'd11027: data <= 8'hFF;
            15'd11028: data <= 8'hFF;
            15'd11029: data <= 8'hFF;
            15'd11030: data <= 8'hFF;
            15'd11031: data <= 8'hFF;
            15'd11032: data <= 8'hFF;
            15'd11033: data <= 8'hFF;
            15'd11034: data <= 8'h80;
            15'd11035: data <= 8'h00;
            15'd11036: data <= 8'h00;
            15'd11037: data <= 8'h00;
            15'd11038: data <= 8'h00;
            15'd11039: data <= 8'h00;
            15'd11040: data <= 8'h00;
            15'd11041: data <= 8'h00;
            15'd11042: data <= 8'h00;
            15'd11043: data <= 8'h00;
            15'd11044: data <= 8'h00;
            15'd11045: data <= 8'h03;
            15'd11046: data <= 8'hFF;
            15'd11047: data <= 8'hFF;
            15'd11048: data <= 8'hFF;
            15'd11049: data <= 8'hFF;
            15'd11050: data <= 8'hFF;
            15'd11051: data <= 8'hFF;
            15'd11052: data <= 8'hFF;
            15'd11053: data <= 8'hFF;
            15'd11054: data <= 8'hFF;
            15'd11055: data <= 8'hFF;
            15'd11056: data <= 8'hFF;
            15'd11057: data <= 8'hFF;
            15'd11058: data <= 8'hFF;
            15'd11059: data <= 8'hFF;
            15'd11060: data <= 8'hFF;
            15'd11061: data <= 8'hFF;
            15'd11062: data <= 8'hFF;
            15'd11063: data <= 8'hFF;
            15'd11064: data <= 8'h80;
            15'd11065: data <= 8'h00;
            15'd11066: data <= 8'h00;
            15'd11067: data <= 8'h00;
            15'd11068: data <= 8'h00;
            15'd11069: data <= 8'h00;
            15'd11070: data <= 8'h00;
            15'd11071: data <= 8'h00;
            15'd11072: data <= 8'h00;
            15'd11073: data <= 8'h00;
            15'd11074: data <= 8'h00;
            15'd11075: data <= 8'h03;
            15'd11076: data <= 8'hFF;
            15'd11077: data <= 8'hFF;
            15'd11078: data <= 8'hFF;
            15'd11079: data <= 8'hFF;
            15'd11080: data <= 8'hFF;
            15'd11081: data <= 8'hFF;
            15'd11082: data <= 8'hFF;
            15'd11083: data <= 8'hFF;
            15'd11084: data <= 8'hFF;
            15'd11085: data <= 8'hFF;
            15'd11086: data <= 8'hFF;
            15'd11087: data <= 8'hFF;
            15'd11088: data <= 8'hFF;
            15'd11089: data <= 8'hFF;
            15'd11090: data <= 8'hFF;
            15'd11091: data <= 8'hFF;
            15'd11092: data <= 8'hFF;
            15'd11093: data <= 8'hFF;
            15'd11094: data <= 8'h80;
            15'd11095: data <= 8'h00;
            15'd11096: data <= 8'h00;
            15'd11097: data <= 8'h00;
            15'd11098: data <= 8'h00;
            15'd11099: data <= 8'h00;
            15'd11100: data <= 8'h00;
            15'd11101: data <= 8'h00;
            15'd11102: data <= 8'h00;
            15'd11103: data <= 8'h00;
            15'd11104: data <= 8'h00;
            15'd11105: data <= 8'h03;
            15'd11106: data <= 8'hFF;
            15'd11107: data <= 8'hFF;
            15'd11108: data <= 8'hFF;
            15'd11109: data <= 8'hFF;
            15'd11110: data <= 8'hFF;
            15'd11111: data <= 8'hFF;
            15'd11112: data <= 8'hFF;
            15'd11113: data <= 8'hFF;
            15'd11114: data <= 8'hFF;
            15'd11115: data <= 8'hFF;
            15'd11116: data <= 8'hFF;
            15'd11117: data <= 8'hFF;
            15'd11118: data <= 8'hFF;
            15'd11119: data <= 8'hFF;
            15'd11120: data <= 8'hFF;
            15'd11121: data <= 8'hFF;
            15'd11122: data <= 8'hFF;
            15'd11123: data <= 8'hFF;
            15'd11124: data <= 8'h80;
            15'd11125: data <= 8'h00;
            15'd11126: data <= 8'h00;
            15'd11127: data <= 8'h00;
            15'd11128: data <= 8'h00;
            15'd11129: data <= 8'h00;
            15'd11130: data <= 8'h00;
            15'd11131: data <= 8'h00;
            15'd11132: data <= 8'h00;
            15'd11133: data <= 8'h00;
            15'd11134: data <= 8'h00;
            15'd11135: data <= 8'h03;
            15'd11136: data <= 8'hFF;
            15'd11137: data <= 8'hFF;
            15'd11138: data <= 8'hFF;
            15'd11139: data <= 8'hFF;
            15'd11140: data <= 8'hFF;
            15'd11141: data <= 8'hFF;
            15'd11142: data <= 8'hFF;
            15'd11143: data <= 8'hFF;
            15'd11144: data <= 8'hFF;
            15'd11145: data <= 8'hFF;
            15'd11146: data <= 8'hFF;
            15'd11147: data <= 8'hFF;
            15'd11148: data <= 8'hFF;
            15'd11149: data <= 8'hFF;
            15'd11150: data <= 8'hFF;
            15'd11151: data <= 8'hFF;
            15'd11152: data <= 8'hFF;
            15'd11153: data <= 8'hFF;
            15'd11154: data <= 8'h80;
            15'd11155: data <= 8'h00;
            15'd11156: data <= 8'h00;
            15'd11157: data <= 8'h00;
            15'd11158: data <= 8'h00;
            15'd11159: data <= 8'h00;
            15'd11160: data <= 8'h00;
            15'd11161: data <= 8'h00;
            15'd11162: data <= 8'h00;
            15'd11163: data <= 8'h00;
            15'd11164: data <= 8'h00;
            15'd11165: data <= 8'h03;
            15'd11166: data <= 8'hFF;
            15'd11167: data <= 8'hFF;
            15'd11168: data <= 8'hFF;
            15'd11169: data <= 8'hFF;
            15'd11170: data <= 8'hFF;
            15'd11171: data <= 8'hFF;
            15'd11172: data <= 8'hFF;
            15'd11173: data <= 8'hFF;
            15'd11174: data <= 8'hFF;
            15'd11175: data <= 8'hFF;
            15'd11176: data <= 8'hFF;
            15'd11177: data <= 8'hFF;
            15'd11178: data <= 8'hFF;
            15'd11179: data <= 8'hFF;
            15'd11180: data <= 8'hFF;
            15'd11181: data <= 8'hFF;
            15'd11182: data <= 8'hFF;
            15'd11183: data <= 8'hFF;
            15'd11184: data <= 8'h80;
            15'd11185: data <= 8'h00;
            15'd11186: data <= 8'h00;
            15'd11187: data <= 8'h00;
            15'd11188: data <= 8'h00;
            15'd11189: data <= 8'h00;
            15'd11190: data <= 8'h00;
            15'd11191: data <= 8'h00;
            15'd11192: data <= 8'h00;
            15'd11193: data <= 8'h00;
            15'd11194: data <= 8'h00;
            15'd11195: data <= 8'h03;
            15'd11196: data <= 8'hFF;
            15'd11197: data <= 8'hFF;
            15'd11198: data <= 8'hFF;
            15'd11199: data <= 8'hFF;
            15'd11200: data <= 8'hFF;
            15'd11201: data <= 8'hFF;
            15'd11202: data <= 8'hFF;
            15'd11203: data <= 8'hFF;
            15'd11204: data <= 8'hFF;
            15'd11205: data <= 8'hFF;
            15'd11206: data <= 8'hFF;
            15'd11207: data <= 8'hFF;
            15'd11208: data <= 8'hFF;
            15'd11209: data <= 8'hFF;
            15'd11210: data <= 8'hFF;
            15'd11211: data <= 8'hFF;
            15'd11212: data <= 8'hFF;
            15'd11213: data <= 8'hFF;
            15'd11214: data <= 8'h80;
            15'd11215: data <= 8'h00;
            15'd11216: data <= 8'h00;
            15'd11217: data <= 8'h00;
            15'd11218: data <= 8'h00;
            15'd11219: data <= 8'h00;
            15'd11220: data <= 8'h00;
            15'd11221: data <= 8'h00;
            15'd11222: data <= 8'h00;
            15'd11223: data <= 8'h00;
            15'd11224: data <= 8'h00;
            15'd11225: data <= 8'h03;
            15'd11226: data <= 8'hFF;
            15'd11227: data <= 8'hFF;
            15'd11228: data <= 8'hFF;
            15'd11229: data <= 8'hFF;
            15'd11230: data <= 8'hFF;
            15'd11231: data <= 8'hFF;
            15'd11232: data <= 8'hFF;
            15'd11233: data <= 8'hFF;
            15'd11234: data <= 8'hFF;
            15'd11235: data <= 8'hFF;
            15'd11236: data <= 8'hFF;
            15'd11237: data <= 8'hFF;
            15'd11238: data <= 8'hFF;
            15'd11239: data <= 8'hFF;
            15'd11240: data <= 8'hFF;
            15'd11241: data <= 8'hFF;
            15'd11242: data <= 8'hFF;
            15'd11243: data <= 8'hFF;
            15'd11244: data <= 8'h80;
            15'd11245: data <= 8'h00;
            15'd11246: data <= 8'h00;
            15'd11247: data <= 8'h00;
            15'd11248: data <= 8'h00;
            15'd11249: data <= 8'h00;
            15'd11250: data <= 8'h00;
            15'd11251: data <= 8'h00;
            15'd11252: data <= 8'h00;
            15'd11253: data <= 8'h00;
            15'd11254: data <= 8'h00;
            15'd11255: data <= 8'h03;
            15'd11256: data <= 8'hFF;
            15'd11257: data <= 8'hFF;
            15'd11258: data <= 8'hFF;
            15'd11259: data <= 8'hFF;
            15'd11260: data <= 8'hFF;
            15'd11261: data <= 8'hFF;
            15'd11262: data <= 8'hFF;
            15'd11263: data <= 8'hFF;
            15'd11264: data <= 8'hFF;
            15'd11265: data <= 8'hFF;
            15'd11266: data <= 8'hFF;
            15'd11267: data <= 8'hFF;
            15'd11268: data <= 8'hFF;
            15'd11269: data <= 8'hFF;
            15'd11270: data <= 8'hFF;
            15'd11271: data <= 8'hFF;
            15'd11272: data <= 8'hFF;
            15'd11273: data <= 8'hFF;
            15'd11274: data <= 8'h80;
            15'd11275: data <= 8'h00;
            15'd11276: data <= 8'h00;
            15'd11277: data <= 8'h00;
            15'd11278: data <= 8'h00;
            15'd11279: data <= 8'h00;
            15'd11280: data <= 8'h00;
            15'd11281: data <= 8'h00;
            15'd11282: data <= 8'h00;
            15'd11283: data <= 8'h00;
            15'd11284: data <= 8'h00;
            15'd11285: data <= 8'h03;
            15'd11286: data <= 8'hFF;
            15'd11287: data <= 8'hFF;
            15'd11288: data <= 8'hFF;
            15'd11289: data <= 8'hFF;
            15'd11290: data <= 8'hFF;
            15'd11291: data <= 8'hFF;
            15'd11292: data <= 8'hFF;
            15'd11293: data <= 8'hFF;
            15'd11294: data <= 8'hFF;
            15'd11295: data <= 8'hFF;
            15'd11296: data <= 8'hFF;
            15'd11297: data <= 8'hFF;
            15'd11298: data <= 8'hFF;
            15'd11299: data <= 8'hFF;
            15'd11300: data <= 8'hFF;
            15'd11301: data <= 8'hFF;
            15'd11302: data <= 8'hFF;
            15'd11303: data <= 8'hFF;
            15'd11304: data <= 8'h80;
            15'd11305: data <= 8'h00;
            15'd11306: data <= 8'h00;
            15'd11307: data <= 8'h00;
            15'd11308: data <= 8'h00;
            15'd11309: data <= 8'h00;
            15'd11310: data <= 8'h00;
            15'd11311: data <= 8'h00;
            15'd11312: data <= 8'h00;
            15'd11313: data <= 8'h00;
            15'd11314: data <= 8'h00;
            15'd11315: data <= 8'h03;
            15'd11316: data <= 8'hFF;
            15'd11317: data <= 8'hFF;
            15'd11318: data <= 8'hFF;
            15'd11319: data <= 8'hFF;
            15'd11320: data <= 8'hFF;
            15'd11321: data <= 8'hFF;
            15'd11322: data <= 8'hFF;
            15'd11323: data <= 8'hFF;
            15'd11324: data <= 8'hFF;
            15'd11325: data <= 8'hFF;
            15'd11326: data <= 8'hFF;
            15'd11327: data <= 8'hFF;
            15'd11328: data <= 8'hFF;
            15'd11329: data <= 8'hFF;
            15'd11330: data <= 8'hFF;
            15'd11331: data <= 8'hFF;
            15'd11332: data <= 8'hFF;
            15'd11333: data <= 8'hFF;
            15'd11334: data <= 8'h80;
            15'd11335: data <= 8'h00;
            15'd11336: data <= 8'h00;
            15'd11337: data <= 8'h00;
            15'd11338: data <= 8'h00;
            15'd11339: data <= 8'h00;
            15'd11340: data <= 8'h00;
            15'd11341: data <= 8'h00;
            15'd11342: data <= 8'h00;
            15'd11343: data <= 8'h00;
            15'd11344: data <= 8'h00;
            15'd11345: data <= 8'h03;
            15'd11346: data <= 8'hFF;
            15'd11347: data <= 8'hFF;
            15'd11348: data <= 8'hFF;
            15'd11349: data <= 8'hFF;
            15'd11350: data <= 8'hFF;
            15'd11351: data <= 8'hFF;
            15'd11352: data <= 8'hFF;
            15'd11353: data <= 8'hFF;
            15'd11354: data <= 8'hFF;
            15'd11355: data <= 8'hFF;
            15'd11356: data <= 8'hFF;
            15'd11357: data <= 8'hFF;
            15'd11358: data <= 8'hFF;
            15'd11359: data <= 8'hFF;
            15'd11360: data <= 8'hFF;
            15'd11361: data <= 8'hFF;
            15'd11362: data <= 8'hFF;
            15'd11363: data <= 8'hFF;
            15'd11364: data <= 8'h80;
            15'd11365: data <= 8'h00;
            15'd11366: data <= 8'h00;
            15'd11367: data <= 8'h00;
            15'd11368: data <= 8'h00;
            15'd11369: data <= 8'h00;
            15'd11370: data <= 8'h00;
            15'd11371: data <= 8'h00;
            15'd11372: data <= 8'h00;
            15'd11373: data <= 8'h00;
            15'd11374: data <= 8'h00;
            15'd11375: data <= 8'h03;
            15'd11376: data <= 8'hFF;
            15'd11377: data <= 8'hFF;
            15'd11378: data <= 8'hFF;
            15'd11379: data <= 8'hFF;
            15'd11380: data <= 8'hFF;
            15'd11381: data <= 8'hFF;
            15'd11382: data <= 8'hFF;
            15'd11383: data <= 8'hFF;
            15'd11384: data <= 8'hFF;
            15'd11385: data <= 8'hFF;
            15'd11386: data <= 8'hFF;
            15'd11387: data <= 8'hFF;
            15'd11388: data <= 8'hFF;
            15'd11389: data <= 8'hFF;
            15'd11390: data <= 8'hFF;
            15'd11391: data <= 8'hFF;
            15'd11392: data <= 8'hFF;
            15'd11393: data <= 8'hFF;
            15'd11394: data <= 8'h80;
            15'd11395: data <= 8'h00;
            15'd11396: data <= 8'h00;
            15'd11397: data <= 8'h00;
            15'd11398: data <= 8'h00;
            15'd11399: data <= 8'h00;
            15'd11400: data <= 8'h00;
            15'd11401: data <= 8'h00;
            15'd11402: data <= 8'h00;
            15'd11403: data <= 8'h00;
            15'd11404: data <= 8'h00;
            15'd11405: data <= 8'h03;
            15'd11406: data <= 8'hFF;
            15'd11407: data <= 8'hFF;
            15'd11408: data <= 8'hFF;
            15'd11409: data <= 8'hFF;
            15'd11410: data <= 8'hFF;
            15'd11411: data <= 8'hFF;
            15'd11412: data <= 8'hFF;
            15'd11413: data <= 8'hFF;
            15'd11414: data <= 8'hFF;
            15'd11415: data <= 8'hFF;
            15'd11416: data <= 8'hFF;
            15'd11417: data <= 8'hFF;
            15'd11418: data <= 8'hFF;
            15'd11419: data <= 8'hFF;
            15'd11420: data <= 8'hFF;
            15'd11421: data <= 8'hFF;
            15'd11422: data <= 8'hFF;
            15'd11423: data <= 8'hFF;
            15'd11424: data <= 8'h80;
            15'd11425: data <= 8'h00;
            15'd11426: data <= 8'h00;
            15'd11427: data <= 8'h00;
            15'd11428: data <= 8'h00;
            15'd11429: data <= 8'h00;
            15'd11430: data <= 8'h00;
            15'd11431: data <= 8'h00;
            15'd11432: data <= 8'h00;
            15'd11433: data <= 8'h00;
            15'd11434: data <= 8'h00;
            15'd11435: data <= 8'h03;
            15'd11436: data <= 8'hFF;
            15'd11437: data <= 8'hFF;
            15'd11438: data <= 8'hFF;
            15'd11439: data <= 8'hFF;
            15'd11440: data <= 8'hFF;
            15'd11441: data <= 8'hFF;
            15'd11442: data <= 8'hFF;
            15'd11443: data <= 8'hFF;
            15'd11444: data <= 8'hFF;
            15'd11445: data <= 8'hFF;
            15'd11446: data <= 8'hFF;
            15'd11447: data <= 8'hFF;
            15'd11448: data <= 8'hFF;
            15'd11449: data <= 8'hFF;
            15'd11450: data <= 8'hFF;
            15'd11451: data <= 8'hFF;
            15'd11452: data <= 8'hFF;
            15'd11453: data <= 8'hFF;
            15'd11454: data <= 8'h80;
            15'd11455: data <= 8'h00;
            15'd11456: data <= 8'h00;
            15'd11457: data <= 8'h00;
            15'd11458: data <= 8'h00;
            15'd11459: data <= 8'h00;
            15'd11460: data <= 8'h00;
            15'd11461: data <= 8'h00;
            15'd11462: data <= 8'h00;
            15'd11463: data <= 8'h00;
            15'd11464: data <= 8'h00;
            15'd11465: data <= 8'h03;
            15'd11466: data <= 8'hFF;
            15'd11467: data <= 8'hFF;
            15'd11468: data <= 8'hFF;
            15'd11469: data <= 8'hFF;
            15'd11470: data <= 8'hFF;
            15'd11471: data <= 8'hFF;
            15'd11472: data <= 8'hFF;
            15'd11473: data <= 8'hFF;
            15'd11474: data <= 8'hFF;
            15'd11475: data <= 8'hFF;
            15'd11476: data <= 8'hFF;
            15'd11477: data <= 8'hFF;
            15'd11478: data <= 8'hFF;
            15'd11479: data <= 8'hFF;
            15'd11480: data <= 8'hFF;
            15'd11481: data <= 8'hFF;
            15'd11482: data <= 8'hFF;
            15'd11483: data <= 8'hFF;
            15'd11484: data <= 8'h80;
            15'd11485: data <= 8'h00;
            15'd11486: data <= 8'h00;
            15'd11487: data <= 8'h00;
            15'd11488: data <= 8'h00;
            15'd11489: data <= 8'h00;
            15'd11490: data <= 8'h00;
            15'd11491: data <= 8'h00;
            15'd11492: data <= 8'h00;
            15'd11493: data <= 8'h00;
            15'd11494: data <= 8'h00;
            15'd11495: data <= 8'h03;
            15'd11496: data <= 8'hFF;
            15'd11497: data <= 8'hFF;
            15'd11498: data <= 8'hFF;
            15'd11499: data <= 8'hFF;
            15'd11500: data <= 8'hFF;
            15'd11501: data <= 8'hFF;
            15'd11502: data <= 8'hFF;
            15'd11503: data <= 8'hFF;
            15'd11504: data <= 8'hFF;
            15'd11505: data <= 8'hFF;
            15'd11506: data <= 8'hFF;
            15'd11507: data <= 8'hFF;
            15'd11508: data <= 8'hFF;
            15'd11509: data <= 8'hFF;
            15'd11510: data <= 8'hFF;
            15'd11511: data <= 8'hFF;
            15'd11512: data <= 8'hFF;
            15'd11513: data <= 8'hFF;
            15'd11514: data <= 8'h80;
            15'd11515: data <= 8'h00;
            15'd11516: data <= 8'h00;
            15'd11517: data <= 8'h00;
            15'd11518: data <= 8'h00;
            15'd11519: data <= 8'h00;
            15'd11520: data <= 8'h00;
            15'd11521: data <= 8'h00;
            15'd11522: data <= 8'h00;
            15'd11523: data <= 8'h00;
            15'd11524: data <= 8'h00;
            15'd11525: data <= 8'h03;
            15'd11526: data <= 8'hFF;
            15'd11527: data <= 8'hFF;
            15'd11528: data <= 8'hFF;
            15'd11529: data <= 8'hFF;
            15'd11530: data <= 8'hFF;
            15'd11531: data <= 8'hFF;
            15'd11532: data <= 8'hFF;
            15'd11533: data <= 8'hFF;
            15'd11534: data <= 8'hFF;
            15'd11535: data <= 8'hFF;
            15'd11536: data <= 8'hFF;
            15'd11537: data <= 8'hFF;
            15'd11538: data <= 8'hFF;
            15'd11539: data <= 8'hFF;
            15'd11540: data <= 8'hFF;
            15'd11541: data <= 8'hFF;
            15'd11542: data <= 8'hFF;
            15'd11543: data <= 8'hFF;
            15'd11544: data <= 8'h80;
            15'd11545: data <= 8'h00;
            15'd11546: data <= 8'h00;
            15'd11547: data <= 8'h00;
            15'd11548: data <= 8'h00;
            15'd11549: data <= 8'h00;
            15'd11550: data <= 8'h00;
            15'd11551: data <= 8'h00;
            15'd11552: data <= 8'h00;
            15'd11553: data <= 8'h00;
            15'd11554: data <= 8'h00;
            15'd11555: data <= 8'h03;
            15'd11556: data <= 8'hFF;
            15'd11557: data <= 8'hFF;
            15'd11558: data <= 8'hFF;
            15'd11559: data <= 8'hFF;
            15'd11560: data <= 8'hFF;
            15'd11561: data <= 8'hFF;
            15'd11562: data <= 8'hFF;
            15'd11563: data <= 8'hFF;
            15'd11564: data <= 8'hFF;
            15'd11565: data <= 8'hFF;
            15'd11566: data <= 8'hFF;
            15'd11567: data <= 8'hFF;
            15'd11568: data <= 8'hFF;
            15'd11569: data <= 8'hFF;
            15'd11570: data <= 8'hFF;
            15'd11571: data <= 8'hFF;
            15'd11572: data <= 8'hFF;
            15'd11573: data <= 8'hFF;
            15'd11574: data <= 8'h80;
            15'd11575: data <= 8'h00;
            15'd11576: data <= 8'h00;
            15'd11577: data <= 8'h00;
            15'd11578: data <= 8'h00;
            15'd11579: data <= 8'h00;
            15'd11580: data <= 8'h00;
            15'd11581: data <= 8'h00;
            15'd11582: data <= 8'h00;
            15'd11583: data <= 8'h00;
            15'd11584: data <= 8'h00;
            15'd11585: data <= 8'h03;
            15'd11586: data <= 8'hFF;
            15'd11587: data <= 8'hFF;
            15'd11588: data <= 8'hFF;
            15'd11589: data <= 8'hFF;
            15'd11590: data <= 8'hFF;
            15'd11591: data <= 8'hFF;
            15'd11592: data <= 8'hFF;
            15'd11593: data <= 8'hFF;
            15'd11594: data <= 8'hFF;
            15'd11595: data <= 8'hFF;
            15'd11596: data <= 8'hFF;
            15'd11597: data <= 8'hFF;
            15'd11598: data <= 8'hFF;
            15'd11599: data <= 8'hFF;
            15'd11600: data <= 8'hFF;
            15'd11601: data <= 8'hFF;
            15'd11602: data <= 8'hFF;
            15'd11603: data <= 8'hFF;
            15'd11604: data <= 8'h80;
            15'd11605: data <= 8'h00;
            15'd11606: data <= 8'h00;
            15'd11607: data <= 8'h00;
            15'd11608: data <= 8'h00;
            15'd11609: data <= 8'h00;
            15'd11610: data <= 8'h00;
            15'd11611: data <= 8'h00;
            15'd11612: data <= 8'h00;
            15'd11613: data <= 8'h00;
            15'd11614: data <= 8'h00;
            15'd11615: data <= 8'h03;
            15'd11616: data <= 8'hFF;
            15'd11617: data <= 8'hFF;
            15'd11618: data <= 8'hFF;
            15'd11619: data <= 8'hFF;
            15'd11620: data <= 8'hFF;
            15'd11621: data <= 8'hFF;
            15'd11622: data <= 8'hFF;
            15'd11623: data <= 8'hFF;
            15'd11624: data <= 8'hFF;
            15'd11625: data <= 8'hFF;
            15'd11626: data <= 8'hFF;
            15'd11627: data <= 8'hFF;
            15'd11628: data <= 8'hFF;
            15'd11629: data <= 8'hFF;
            15'd11630: data <= 8'hFF;
            15'd11631: data <= 8'hFF;
            15'd11632: data <= 8'hFF;
            15'd11633: data <= 8'hFF;
            15'd11634: data <= 8'h80;
            15'd11635: data <= 8'h00;
            15'd11636: data <= 8'h00;
            15'd11637: data <= 8'h00;
            15'd11638: data <= 8'h00;
            15'd11639: data <= 8'h00;
            15'd11640: data <= 8'h00;
            15'd11641: data <= 8'h00;
            15'd11642: data <= 8'h00;
            15'd11643: data <= 8'h00;
            15'd11644: data <= 8'h00;
            15'd11645: data <= 8'h03;
            15'd11646: data <= 8'hFF;
            15'd11647: data <= 8'hFF;
            15'd11648: data <= 8'hFF;
            15'd11649: data <= 8'hFF;
            15'd11650: data <= 8'hFF;
            15'd11651: data <= 8'hFF;
            15'd11652: data <= 8'hFF;
            15'd11653: data <= 8'hFF;
            15'd11654: data <= 8'hFF;
            15'd11655: data <= 8'hFF;
            15'd11656: data <= 8'hFF;
            15'd11657: data <= 8'hFF;
            15'd11658: data <= 8'hFF;
            15'd11659: data <= 8'hFF;
            15'd11660: data <= 8'hFF;
            15'd11661: data <= 8'hFF;
            15'd11662: data <= 8'hFF;
            15'd11663: data <= 8'hFF;
            15'd11664: data <= 8'h80;
            15'd11665: data <= 8'h00;
            15'd11666: data <= 8'h00;
            15'd11667: data <= 8'h00;
            15'd11668: data <= 8'h00;
            15'd11669: data <= 8'h00;
            15'd11670: data <= 8'h00;
            15'd11671: data <= 8'h00;
            15'd11672: data <= 8'h00;
            15'd11673: data <= 8'h00;
            15'd11674: data <= 8'h00;
            15'd11675: data <= 8'h03;
            15'd11676: data <= 8'hFF;
            15'd11677: data <= 8'hFF;
            15'd11678: data <= 8'hFF;
            15'd11679: data <= 8'hFF;
            15'd11680: data <= 8'hFF;
            15'd11681: data <= 8'hFF;
            15'd11682: data <= 8'hFF;
            15'd11683: data <= 8'hFF;
            15'd11684: data <= 8'hFF;
            15'd11685: data <= 8'hFF;
            15'd11686: data <= 8'hFF;
            15'd11687: data <= 8'hFF;
            15'd11688: data <= 8'hFF;
            15'd11689: data <= 8'hFF;
            15'd11690: data <= 8'hFF;
            15'd11691: data <= 8'hFF;
            15'd11692: data <= 8'hFF;
            15'd11693: data <= 8'hFF;
            15'd11694: data <= 8'h80;
            15'd11695: data <= 8'h00;
            15'd11696: data <= 8'h00;
            15'd11697: data <= 8'h00;
            15'd11698: data <= 8'h00;
            15'd11699: data <= 8'h00;
            15'd11700: data <= 8'h00;
            15'd11701: data <= 8'h00;
            15'd11702: data <= 8'h00;
            15'd11703: data <= 8'h00;
            15'd11704: data <= 8'h00;
            15'd11705: data <= 8'h03;
            15'd11706: data <= 8'hFF;
            15'd11707: data <= 8'hFF;
            15'd11708: data <= 8'hFF;
            15'd11709: data <= 8'hFF;
            15'd11710: data <= 8'hFF;
            15'd11711: data <= 8'hFF;
            15'd11712: data <= 8'hFF;
            15'd11713: data <= 8'hFF;
            15'd11714: data <= 8'hFF;
            15'd11715: data <= 8'hE0;
            15'd11716: data <= 8'hFF;
            15'd11717: data <= 8'hFF;
            15'd11718: data <= 8'hFF;
            15'd11719: data <= 8'hFF;
            15'd11720: data <= 8'hFF;
            15'd11721: data <= 8'hFF;
            15'd11722: data <= 8'hFF;
            15'd11723: data <= 8'hFF;
            15'd11724: data <= 8'h80;
            15'd11725: data <= 8'h00;
            15'd11726: data <= 8'h00;
            15'd11727: data <= 8'h00;
            15'd11728: data <= 8'h00;
            15'd11729: data <= 8'h00;
            15'd11730: data <= 8'h00;
            15'd11731: data <= 8'h00;
            15'd11732: data <= 8'h00;
            15'd11733: data <= 8'h00;
            15'd11734: data <= 8'h00;
            15'd11735: data <= 8'h03;
            15'd11736: data <= 8'hFF;
            15'd11737: data <= 8'hFF;
            15'd11738: data <= 8'hFF;
            15'd11739: data <= 8'hFF;
            15'd11740: data <= 8'hFF;
            15'd11741: data <= 8'hFF;
            15'd11742: data <= 8'hFF;
            15'd11743: data <= 8'hFF;
            15'd11744: data <= 8'hFF;
            15'd11745: data <= 8'h80;
            15'd11746: data <= 8'h3F;
            15'd11747: data <= 8'hFF;
            15'd11748: data <= 8'hFF;
            15'd11749: data <= 8'hFF;
            15'd11750: data <= 8'hFF;
            15'd11751: data <= 8'hFF;
            15'd11752: data <= 8'hFF;
            15'd11753: data <= 8'hFF;
            15'd11754: data <= 8'h80;
            15'd11755: data <= 8'h00;
            15'd11756: data <= 8'h00;
            15'd11757: data <= 8'h00;
            15'd11758: data <= 8'h00;
            15'd11759: data <= 8'h00;
            15'd11760: data <= 8'h00;
            15'd11761: data <= 8'h00;
            15'd11762: data <= 8'h00;
            15'd11763: data <= 8'h00;
            15'd11764: data <= 8'h00;
            15'd11765: data <= 8'h03;
            15'd11766: data <= 8'hFF;
            15'd11767: data <= 8'hFF;
            15'd11768: data <= 8'hFF;
            15'd11769: data <= 8'hFF;
            15'd11770: data <= 8'hFF;
            15'd11771: data <= 8'hFF;
            15'd11772: data <= 8'hFF;
            15'd11773: data <= 8'hFF;
            15'd11774: data <= 8'h80;
            15'd11775: data <= 8'h00;
            15'd11776: data <= 8'h1F;
            15'd11777: data <= 8'hFF;
            15'd11778: data <= 8'hFF;
            15'd11779: data <= 8'hFF;
            15'd11780: data <= 8'hFF;
            15'd11781: data <= 8'hFF;
            15'd11782: data <= 8'hFF;
            15'd11783: data <= 8'hFF;
            15'd11784: data <= 8'h80;
            15'd11785: data <= 8'h00;
            15'd11786: data <= 8'h00;
            15'd11787: data <= 8'h00;
            15'd11788: data <= 8'h00;
            15'd11789: data <= 8'h00;
            15'd11790: data <= 8'h00;
            15'd11791: data <= 8'h00;
            15'd11792: data <= 8'h00;
            15'd11793: data <= 8'h00;
            15'd11794: data <= 8'h00;
            15'd11795: data <= 8'h03;
            15'd11796: data <= 8'hFF;
            15'd11797: data <= 8'hFF;
            15'd11798: data <= 8'hFF;
            15'd11799: data <= 8'hFF;
            15'd11800: data <= 8'hFF;
            15'd11801: data <= 8'hFF;
            15'd11802: data <= 8'hFF;
            15'd11803: data <= 8'h80;
            15'd11804: data <= 8'h00;
            15'd11805: data <= 8'h00;
            15'd11806: data <= 8'h1F;
            15'd11807: data <= 8'hFF;
            15'd11808: data <= 8'hFF;
            15'd11809: data <= 8'hFF;
            15'd11810: data <= 8'hFF;
            15'd11811: data <= 8'hFF;
            15'd11812: data <= 8'hFF;
            15'd11813: data <= 8'hFF;
            15'd11814: data <= 8'h80;
            15'd11815: data <= 8'h00;
            15'd11816: data <= 8'h00;
            15'd11817: data <= 8'h00;
            15'd11818: data <= 8'h00;
            15'd11819: data <= 8'h00;
            15'd11820: data <= 8'h00;
            15'd11821: data <= 8'h00;
            15'd11822: data <= 8'h00;
            15'd11823: data <= 8'h00;
            15'd11824: data <= 8'h00;
            15'd11825: data <= 8'h03;
            15'd11826: data <= 8'hFF;
            15'd11827: data <= 8'hFF;
            15'd11828: data <= 8'hFF;
            15'd11829: data <= 8'hFF;
            15'd11830: data <= 8'hFF;
            15'd11831: data <= 8'hFF;
            15'd11832: data <= 8'hFE;
            15'd11833: data <= 8'h00;
            15'd11834: data <= 8'h00;
            15'd11835: data <= 8'h00;
            15'd11836: data <= 8'h1F;
            15'd11837: data <= 8'hFF;
            15'd11838: data <= 8'hFF;
            15'd11839: data <= 8'hFF;
            15'd11840: data <= 8'hFF;
            15'd11841: data <= 8'hFF;
            15'd11842: data <= 8'hFF;
            15'd11843: data <= 8'hFF;
            15'd11844: data <= 8'h80;
            15'd11845: data <= 8'h00;
            15'd11846: data <= 8'h00;
            15'd11847: data <= 8'h00;
            15'd11848: data <= 8'h00;
            15'd11849: data <= 8'h00;
            15'd11850: data <= 8'h00;
            15'd11851: data <= 8'h00;
            15'd11852: data <= 8'h00;
            15'd11853: data <= 8'h00;
            15'd11854: data <= 8'h00;
            15'd11855: data <= 8'h03;
            15'd11856: data <= 8'hFF;
            15'd11857: data <= 8'hFF;
            15'd11858: data <= 8'hFF;
            15'd11859: data <= 8'hFF;
            15'd11860: data <= 8'hFF;
            15'd11861: data <= 8'hFF;
            15'd11862: data <= 8'h80;
            15'd11863: data <= 8'h00;
            15'd11864: data <= 8'h00;
            15'd11865: data <= 8'h00;
            15'd11866: data <= 8'h0F;
            15'd11867: data <= 8'hFF;
            15'd11868: data <= 8'hFF;
            15'd11869: data <= 8'hFF;
            15'd11870: data <= 8'hFF;
            15'd11871: data <= 8'hFF;
            15'd11872: data <= 8'hFF;
            15'd11873: data <= 8'hFF;
            15'd11874: data <= 8'h80;
            15'd11875: data <= 8'h00;
            15'd11876: data <= 8'h00;
            15'd11877: data <= 8'h00;
            15'd11878: data <= 8'h00;
            15'd11879: data <= 8'h00;
            15'd11880: data <= 8'h00;
            15'd11881: data <= 8'h00;
            15'd11882: data <= 8'h00;
            15'd11883: data <= 8'h00;
            15'd11884: data <= 8'h00;
            15'd11885: data <= 8'h03;
            15'd11886: data <= 8'hFF;
            15'd11887: data <= 8'hFF;
            15'd11888: data <= 8'hFF;
            15'd11889: data <= 8'hFF;
            15'd11890: data <= 8'hFF;
            15'd11891: data <= 8'hFE;
            15'd11892: data <= 8'h00;
            15'd11893: data <= 8'h00;
            15'd11894: data <= 8'h00;
            15'd11895: data <= 8'h00;
            15'd11896: data <= 8'h07;
            15'd11897: data <= 8'hFF;
            15'd11898: data <= 8'hFF;
            15'd11899: data <= 8'hFF;
            15'd11900: data <= 8'hFF;
            15'd11901: data <= 8'hFF;
            15'd11902: data <= 8'hFF;
            15'd11903: data <= 8'hFF;
            15'd11904: data <= 8'h80;
            15'd11905: data <= 8'h00;
            15'd11906: data <= 8'h00;
            15'd11907: data <= 8'h00;
            15'd11908: data <= 8'h00;
            15'd11909: data <= 8'h00;
            15'd11910: data <= 8'h00;
            15'd11911: data <= 8'h00;
            15'd11912: data <= 8'h00;
            15'd11913: data <= 8'h00;
            15'd11914: data <= 8'h00;
            15'd11915: data <= 8'h03;
            15'd11916: data <= 8'hFF;
            15'd11917: data <= 8'hFF;
            15'd11918: data <= 8'hFF;
            15'd11919: data <= 8'hFF;
            15'd11920: data <= 8'hFF;
            15'd11921: data <= 8'hF0;
            15'd11922: data <= 8'h00;
            15'd11923: data <= 8'h00;
            15'd11924: data <= 8'h00;
            15'd11925: data <= 8'h10;
            15'd11926: data <= 8'h07;
            15'd11927: data <= 8'hFF;
            15'd11928: data <= 8'hFF;
            15'd11929: data <= 8'hFF;
            15'd11930: data <= 8'hFF;
            15'd11931: data <= 8'hFF;
            15'd11932: data <= 8'hFF;
            15'd11933: data <= 8'hFF;
            15'd11934: data <= 8'h80;
            15'd11935: data <= 8'h00;
            15'd11936: data <= 8'h00;
            15'd11937: data <= 8'h00;
            15'd11938: data <= 8'h00;
            15'd11939: data <= 8'h00;
            15'd11940: data <= 8'h00;
            15'd11941: data <= 8'h00;
            15'd11942: data <= 8'h00;
            15'd11943: data <= 8'h00;
            15'd11944: data <= 8'h00;
            15'd11945: data <= 8'h03;
            15'd11946: data <= 8'hFF;
            15'd11947: data <= 8'hFF;
            15'd11948: data <= 8'hFF;
            15'd11949: data <= 8'hFF;
            15'd11950: data <= 8'hFF;
            15'd11951: data <= 8'hC0;
            15'd11952: data <= 8'h00;
            15'd11953: data <= 8'h00;
            15'd11954: data <= 8'h01;
            15'd11955: data <= 8'hFC;
            15'd11956: data <= 8'h03;
            15'd11957: data <= 8'hFF;
            15'd11958: data <= 8'hFF;
            15'd11959: data <= 8'hFF;
            15'd11960: data <= 8'hFF;
            15'd11961: data <= 8'hFF;
            15'd11962: data <= 8'hFF;
            15'd11963: data <= 8'hFF;
            15'd11964: data <= 8'h80;
            15'd11965: data <= 8'h00;
            15'd11966: data <= 8'h00;
            15'd11967: data <= 8'h00;
            15'd11968: data <= 8'h00;
            15'd11969: data <= 8'h00;
            15'd11970: data <= 8'h00;
            15'd11971: data <= 8'h00;
            15'd11972: data <= 8'h00;
            15'd11973: data <= 8'h00;
            15'd11974: data <= 8'h00;
            15'd11975: data <= 8'h03;
            15'd11976: data <= 8'hFF;
            15'd11977: data <= 8'hFF;
            15'd11978: data <= 8'hFF;
            15'd11979: data <= 8'hFF;
            15'd11980: data <= 8'hFE;
            15'd11981: data <= 8'h00;
            15'd11982: data <= 8'h00;
            15'd11983: data <= 8'h00;
            15'd11984: data <= 8'hFF;
            15'd11985: data <= 8'hFE;
            15'd11986: data <= 8'h00;
            15'd11987: data <= 8'h7F;
            15'd11988: data <= 8'hFF;
            15'd11989: data <= 8'hFF;
            15'd11990: data <= 8'hFF;
            15'd11991: data <= 8'hFF;
            15'd11992: data <= 8'hFF;
            15'd11993: data <= 8'hFF;
            15'd11994: data <= 8'h80;
            15'd11995: data <= 8'h00;
            15'd11996: data <= 8'h00;
            15'd11997: data <= 8'h00;
            15'd11998: data <= 8'h00;
            15'd11999: data <= 8'h00;
            15'd12000: data <= 8'h00;
            15'd12001: data <= 8'h00;
            15'd12002: data <= 8'h00;
            15'd12003: data <= 8'h00;
            15'd12004: data <= 8'h00;
            15'd12005: data <= 8'h03;
            15'd12006: data <= 8'hFF;
            15'd12007: data <= 8'hFF;
            15'd12008: data <= 8'hFF;
            15'd12009: data <= 8'hFF;
            15'd12010: data <= 8'hF8;
            15'd12011: data <= 8'h00;
            15'd12012: data <= 8'h00;
            15'd12013: data <= 8'h3F;
            15'd12014: data <= 8'hFF;
            15'd12015: data <= 8'hFE;
            15'd12016: data <= 8'h00;
            15'd12017: data <= 8'h1F;
            15'd12018: data <= 8'hFF;
            15'd12019: data <= 8'hFF;
            15'd12020: data <= 8'hFF;
            15'd12021: data <= 8'hFF;
            15'd12022: data <= 8'hFF;
            15'd12023: data <= 8'hFF;
            15'd12024: data <= 8'h80;
            15'd12025: data <= 8'h00;
            15'd12026: data <= 8'h00;
            15'd12027: data <= 8'h00;
            15'd12028: data <= 8'h00;
            15'd12029: data <= 8'h00;
            15'd12030: data <= 8'h00;
            15'd12031: data <= 8'h00;
            15'd12032: data <= 8'h00;
            15'd12033: data <= 8'h00;
            15'd12034: data <= 8'h00;
            15'd12035: data <= 8'h03;
            15'd12036: data <= 8'hFF;
            15'd12037: data <= 8'hFF;
            15'd12038: data <= 8'hFF;
            15'd12039: data <= 8'hFF;
            15'd12040: data <= 8'hC0;
            15'd12041: data <= 8'h00;
            15'd12042: data <= 8'h07;
            15'd12043: data <= 8'hFF;
            15'd12044: data <= 8'hFF;
            15'd12045: data <= 8'hFF;
            15'd12046: data <= 8'h00;
            15'd12047: data <= 8'h03;
            15'd12048: data <= 8'hFF;
            15'd12049: data <= 8'hFF;
            15'd12050: data <= 8'hFF;
            15'd12051: data <= 8'hFF;
            15'd12052: data <= 8'hFF;
            15'd12053: data <= 8'hFF;
            15'd12054: data <= 8'h80;
            15'd12055: data <= 8'h00;
            15'd12056: data <= 8'h00;
            15'd12057: data <= 8'h00;
            15'd12058: data <= 8'h00;
            15'd12059: data <= 8'h00;
            15'd12060: data <= 8'h00;
            15'd12061: data <= 8'h00;
            15'd12062: data <= 8'h00;
            15'd12063: data <= 8'h00;
            15'd12064: data <= 8'h00;
            15'd12065: data <= 8'h03;
            15'd12066: data <= 8'hFF;
            15'd12067: data <= 8'hFF;
            15'd12068: data <= 8'hFF;
            15'd12069: data <= 8'hFF;
            15'd12070: data <= 8'h00;
            15'd12071: data <= 8'h00;
            15'd12072: data <= 8'h3F;
            15'd12073: data <= 8'hFF;
            15'd12074: data <= 8'hFF;
            15'd12075: data <= 8'hFF;
            15'd12076: data <= 8'h80;
            15'd12077: data <= 8'h00;
            15'd12078: data <= 8'h7F;
            15'd12079: data <= 8'hFF;
            15'd12080: data <= 8'hFF;
            15'd12081: data <= 8'hFF;
            15'd12082: data <= 8'hFF;
            15'd12083: data <= 8'hFF;
            15'd12084: data <= 8'h80;
            15'd12085: data <= 8'h00;
            15'd12086: data <= 8'h00;
            15'd12087: data <= 8'h00;
            15'd12088: data <= 8'h00;
            15'd12089: data <= 8'h00;
            15'd12090: data <= 8'h00;
            15'd12091: data <= 8'h00;
            15'd12092: data <= 8'h00;
            15'd12093: data <= 8'h00;
            15'd12094: data <= 8'h00;
            15'd12095: data <= 8'h03;
            15'd12096: data <= 8'hFF;
            15'd12097: data <= 8'hFF;
            15'd12098: data <= 8'hFF;
            15'd12099: data <= 8'hFE;
            15'd12100: data <= 8'h00;
            15'd12101: data <= 8'h01;
            15'd12102: data <= 8'hFF;
            15'd12103: data <= 8'hFF;
            15'd12104: data <= 8'hFF;
            15'd12105: data <= 8'hFF;
            15'd12106: data <= 8'hC0;
            15'd12107: data <= 8'h00;
            15'd12108: data <= 8'h04;
            15'd12109: data <= 8'h03;
            15'd12110: data <= 8'hFF;
            15'd12111: data <= 8'hFF;
            15'd12112: data <= 8'hFF;
            15'd12113: data <= 8'hFF;
            15'd12114: data <= 8'h80;
            15'd12115: data <= 8'h00;
            15'd12116: data <= 8'h00;
            15'd12117: data <= 8'h00;
            15'd12118: data <= 8'h00;
            15'd12119: data <= 8'h00;
            15'd12120: data <= 8'h00;
            15'd12121: data <= 8'h00;
            15'd12122: data <= 8'h00;
            15'd12123: data <= 8'h00;
            15'd12124: data <= 8'h00;
            15'd12125: data <= 8'h03;
            15'd12126: data <= 8'hFF;
            15'd12127: data <= 8'hFF;
            15'd12128: data <= 8'hFF;
            15'd12129: data <= 8'hFC;
            15'd12130: data <= 8'h00;
            15'd12131: data <= 8'h0F;
            15'd12132: data <= 8'hFF;
            15'd12133: data <= 8'hFF;
            15'd12134: data <= 8'hFF;
            15'd12135: data <= 8'hFF;
            15'd12136: data <= 8'hF0;
            15'd12137: data <= 8'h00;
            15'd12138: data <= 8'h00;
            15'd12139: data <= 8'h01;
            15'd12140: data <= 8'hFF;
            15'd12141: data <= 8'hFF;
            15'd12142: data <= 8'hFF;
            15'd12143: data <= 8'hFF;
            15'd12144: data <= 8'h80;
            15'd12145: data <= 8'h00;
            15'd12146: data <= 8'h00;
            15'd12147: data <= 8'h00;
            15'd12148: data <= 8'h00;
            15'd12149: data <= 8'h00;
            15'd12150: data <= 8'h00;
            15'd12151: data <= 8'h00;
            15'd12152: data <= 8'h00;
            15'd12153: data <= 8'h00;
            15'd12154: data <= 8'h00;
            15'd12155: data <= 8'h03;
            15'd12156: data <= 8'hFF;
            15'd12157: data <= 8'hFF;
            15'd12158: data <= 8'hFF;
            15'd12159: data <= 8'hF0;
            15'd12160: data <= 8'h00;
            15'd12161: data <= 8'h7F;
            15'd12162: data <= 8'hFF;
            15'd12163: data <= 8'hFF;
            15'd12164: data <= 8'hFF;
            15'd12165: data <= 8'hFF;
            15'd12166: data <= 8'hFC;
            15'd12167: data <= 8'h00;
            15'd12168: data <= 8'h00;
            15'd12169: data <= 8'h00;
            15'd12170: data <= 8'hFF;
            15'd12171: data <= 8'hFF;
            15'd12172: data <= 8'hFF;
            15'd12173: data <= 8'hFF;
            15'd12174: data <= 8'h80;
            15'd12175: data <= 8'h00;
            15'd12176: data <= 8'h00;
            15'd12177: data <= 8'h00;
            15'd12178: data <= 8'h00;
            15'd12179: data <= 8'h00;
            15'd12180: data <= 8'h00;
            15'd12181: data <= 8'h00;
            15'd12182: data <= 8'h00;
            15'd12183: data <= 8'h00;
            15'd12184: data <= 8'h00;
            15'd12185: data <= 8'h03;
            15'd12186: data <= 8'hFF;
            15'd12187: data <= 8'hFF;
            15'd12188: data <= 8'hFF;
            15'd12189: data <= 8'hE0;
            15'd12190: data <= 8'h03;
            15'd12191: data <= 8'hFF;
            15'd12192: data <= 8'hFF;
            15'd12193: data <= 8'hFF;
            15'd12194: data <= 8'hFF;
            15'd12195: data <= 8'hFF;
            15'd12196: data <= 8'hFF;
            15'd12197: data <= 8'h00;
            15'd12198: data <= 8'h00;
            15'd12199: data <= 8'h00;
            15'd12200: data <= 8'h7F;
            15'd12201: data <= 8'hFF;
            15'd12202: data <= 8'hFF;
            15'd12203: data <= 8'hFF;
            15'd12204: data <= 8'h80;
            15'd12205: data <= 8'h00;
            15'd12206: data <= 8'h00;
            15'd12207: data <= 8'h00;
            15'd12208: data <= 8'h00;
            15'd12209: data <= 8'h00;
            15'd12210: data <= 8'h00;
            15'd12211: data <= 8'h00;
            15'd12212: data <= 8'h00;
            15'd12213: data <= 8'h00;
            15'd12214: data <= 8'h00;
            15'd12215: data <= 8'h03;
            15'd12216: data <= 8'hFF;
            15'd12217: data <= 8'hFF;
            15'd12218: data <= 8'hFF;
            15'd12219: data <= 8'h80;
            15'd12220: data <= 8'h07;
            15'd12221: data <= 8'hFF;
            15'd12222: data <= 8'hFF;
            15'd12223: data <= 8'hFF;
            15'd12224: data <= 8'hFF;
            15'd12225: data <= 8'hFF;
            15'd12226: data <= 8'hFF;
            15'd12227: data <= 8'hE0;
            15'd12228: data <= 8'h00;
            15'd12229: data <= 8'h00;
            15'd12230: data <= 8'h7F;
            15'd12231: data <= 8'hFF;
            15'd12232: data <= 8'hFF;
            15'd12233: data <= 8'hFF;
            15'd12234: data <= 8'h80;
            15'd12235: data <= 8'h00;
            15'd12236: data <= 8'h00;
            15'd12237: data <= 8'h00;
            15'd12238: data <= 8'h00;
            15'd12239: data <= 8'h00;
            15'd12240: data <= 8'h00;
            15'd12241: data <= 8'h00;
            15'd12242: data <= 8'h00;
            15'd12243: data <= 8'h00;
            15'd12244: data <= 8'h00;
            15'd12245: data <= 8'h03;
            15'd12246: data <= 8'hFF;
            15'd12247: data <= 8'hFF;
            15'd12248: data <= 8'hFF;
            15'd12249: data <= 8'h00;
            15'd12250: data <= 8'h0F;
            15'd12251: data <= 8'hFF;
            15'd12252: data <= 8'hFF;
            15'd12253: data <= 8'hFF;
            15'd12254: data <= 8'hFF;
            15'd12255: data <= 8'hFF;
            15'd12256: data <= 8'hFF;
            15'd12257: data <= 8'hFE;
            15'd12258: data <= 8'h00;
            15'd12259: data <= 8'h00;
            15'd12260: data <= 8'h3F;
            15'd12261: data <= 8'hFF;
            15'd12262: data <= 8'hFF;
            15'd12263: data <= 8'hFF;
            15'd12264: data <= 8'h80;
            15'd12265: data <= 8'h00;
            15'd12266: data <= 8'h00;
            15'd12267: data <= 8'h00;
            15'd12268: data <= 8'h00;
            15'd12269: data <= 8'h00;
            15'd12270: data <= 8'h00;
            15'd12271: data <= 8'h00;
            15'd12272: data <= 8'h00;
            15'd12273: data <= 8'h00;
            15'd12274: data <= 8'h00;
            15'd12275: data <= 8'h03;
            15'd12276: data <= 8'hFF;
            15'd12277: data <= 8'hFF;
            15'd12278: data <= 8'hFE;
            15'd12279: data <= 8'h00;
            15'd12280: data <= 8'h3F;
            15'd12281: data <= 8'hFF;
            15'd12282: data <= 8'hFF;
            15'd12283: data <= 8'hFF;
            15'd12284: data <= 8'hFF;
            15'd12285: data <= 8'hFF;
            15'd12286: data <= 8'hFF;
            15'd12287: data <= 8'hFF;
            15'd12288: data <= 8'h80;
            15'd12289: data <= 8'h00;
            15'd12290: data <= 8'h3F;
            15'd12291: data <= 8'hFF;
            15'd12292: data <= 8'hFF;
            15'd12293: data <= 8'hFF;
            15'd12294: data <= 8'h80;
            15'd12295: data <= 8'h00;
            15'd12296: data <= 8'h00;
            15'd12297: data <= 8'h00;
            15'd12298: data <= 8'h00;
            15'd12299: data <= 8'h00;
            15'd12300: data <= 8'h00;
            15'd12301: data <= 8'h00;
            15'd12302: data <= 8'h00;
            15'd12303: data <= 8'h00;
            15'd12304: data <= 8'h00;
            15'd12305: data <= 8'h03;
            15'd12306: data <= 8'hFF;
            15'd12307: data <= 8'hFF;
            15'd12308: data <= 8'hFC;
            15'd12309: data <= 8'h00;
            15'd12310: data <= 8'hFF;
            15'd12311: data <= 8'hFF;
            15'd12312: data <= 8'hFF;
            15'd12313: data <= 8'hFF;
            15'd12314: data <= 8'hFF;
            15'd12315: data <= 8'hFF;
            15'd12316: data <= 8'hFF;
            15'd12317: data <= 8'hFF;
            15'd12318: data <= 8'hFF;
            15'd12319: data <= 8'hE0;
            15'd12320: data <= 8'h3F;
            15'd12321: data <= 8'hFF;
            15'd12322: data <= 8'hFF;
            15'd12323: data <= 8'hFF;
            15'd12324: data <= 8'h80;
            15'd12325: data <= 8'h00;
            15'd12326: data <= 8'h00;
            15'd12327: data <= 8'h00;
            15'd12328: data <= 8'h00;
            15'd12329: data <= 8'h00;
            15'd12330: data <= 8'h00;
            15'd12331: data <= 8'h00;
            15'd12332: data <= 8'h00;
            15'd12333: data <= 8'h00;
            15'd12334: data <= 8'h00;
            15'd12335: data <= 8'h03;
            15'd12336: data <= 8'hFF;
            15'd12337: data <= 8'hFF;
            15'd12338: data <= 8'hF8;
            15'd12339: data <= 8'h01;
            15'd12340: data <= 8'hFF;
            15'd12341: data <= 8'hFF;
            15'd12342: data <= 8'hFF;
            15'd12343: data <= 8'hFF;
            15'd12344: data <= 8'hFF;
            15'd12345: data <= 8'hFF;
            15'd12346: data <= 8'hFF;
            15'd12347: data <= 8'hFF;
            15'd12348: data <= 8'hFF;
            15'd12349: data <= 8'hF0;
            15'd12350: data <= 8'h1F;
            15'd12351: data <= 8'hFF;
            15'd12352: data <= 8'hFF;
            15'd12353: data <= 8'hFF;
            15'd12354: data <= 8'h80;
            15'd12355: data <= 8'h00;
            15'd12356: data <= 8'h00;
            15'd12357: data <= 8'h00;
            15'd12358: data <= 8'h00;
            15'd12359: data <= 8'h00;
            15'd12360: data <= 8'h00;
            15'd12361: data <= 8'h00;
            15'd12362: data <= 8'h00;
            15'd12363: data <= 8'h00;
            15'd12364: data <= 8'h00;
            15'd12365: data <= 8'h03;
            15'd12366: data <= 8'hFF;
            15'd12367: data <= 8'hFF;
            15'd12368: data <= 8'hF0;
            15'd12369: data <= 8'h03;
            15'd12370: data <= 8'hFF;
            15'd12371: data <= 8'hFF;
            15'd12372: data <= 8'hFF;
            15'd12373: data <= 8'hFF;
            15'd12374: data <= 8'hFF;
            15'd12375: data <= 8'hFF;
            15'd12376: data <= 8'hFF;
            15'd12377: data <= 8'hFF;
            15'd12378: data <= 8'hFF;
            15'd12379: data <= 8'hF0;
            15'd12380: data <= 8'h1F;
            15'd12381: data <= 8'hFF;
            15'd12382: data <= 8'hFF;
            15'd12383: data <= 8'hFF;
            15'd12384: data <= 8'h80;
            15'd12385: data <= 8'h00;
            15'd12386: data <= 8'h00;
            15'd12387: data <= 8'h00;
            15'd12388: data <= 8'h00;
            15'd12389: data <= 8'h00;
            15'd12390: data <= 8'h00;
            15'd12391: data <= 8'h00;
            15'd12392: data <= 8'h00;
            15'd12393: data <= 8'h00;
            15'd12394: data <= 8'h00;
            15'd12395: data <= 8'h03;
            15'd12396: data <= 8'hFF;
            15'd12397: data <= 8'hFF;
            15'd12398: data <= 8'hF0;
            15'd12399: data <= 8'h0F;
            15'd12400: data <= 8'hFF;
            15'd12401: data <= 8'hFF;
            15'd12402: data <= 8'hFF;
            15'd12403: data <= 8'hFF;
            15'd12404: data <= 8'hFF;
            15'd12405: data <= 8'hFF;
            15'd12406: data <= 8'hFF;
            15'd12407: data <= 8'hFF;
            15'd12408: data <= 8'hFF;
            15'd12409: data <= 8'hF0;
            15'd12410: data <= 8'h1F;
            15'd12411: data <= 8'hFF;
            15'd12412: data <= 8'hFF;
            15'd12413: data <= 8'hFF;
            15'd12414: data <= 8'h80;
            15'd12415: data <= 8'h00;
            15'd12416: data <= 8'h00;
            15'd12417: data <= 8'h00;
            15'd12418: data <= 8'h00;
            15'd12419: data <= 8'h00;
            15'd12420: data <= 8'h00;
            15'd12421: data <= 8'h00;
            15'd12422: data <= 8'h00;
            15'd12423: data <= 8'h00;
            15'd12424: data <= 8'h00;
            15'd12425: data <= 8'h03;
            15'd12426: data <= 8'hFF;
            15'd12427: data <= 8'hFF;
            15'd12428: data <= 8'hE0;
            15'd12429: data <= 8'h0F;
            15'd12430: data <= 8'hFF;
            15'd12431: data <= 8'hFF;
            15'd12432: data <= 8'hFF;
            15'd12433: data <= 8'hFF;
            15'd12434: data <= 8'hFF;
            15'd12435: data <= 8'hFF;
            15'd12436: data <= 8'hFF;
            15'd12437: data <= 8'hFF;
            15'd12438: data <= 8'hFF;
            15'd12439: data <= 8'hF8;
            15'd12440: data <= 8'h0F;
            15'd12441: data <= 8'hFF;
            15'd12442: data <= 8'hFF;
            15'd12443: data <= 8'hFF;
            15'd12444: data <= 8'h80;
            15'd12445: data <= 8'h00;
            15'd12446: data <= 8'h00;
            15'd12447: data <= 8'h00;
            15'd12448: data <= 8'h00;
            15'd12449: data <= 8'h00;
            15'd12450: data <= 8'h00;
            15'd12451: data <= 8'h00;
            15'd12452: data <= 8'h00;
            15'd12453: data <= 8'h00;
            15'd12454: data <= 8'h00;
            15'd12455: data <= 8'h03;
            15'd12456: data <= 8'hFF;
            15'd12457: data <= 8'hFF;
            15'd12458: data <= 8'hC0;
            15'd12459: data <= 8'h1F;
            15'd12460: data <= 8'hFF;
            15'd12461: data <= 8'hFF;
            15'd12462: data <= 8'hFF;
            15'd12463: data <= 8'hFF;
            15'd12464: data <= 8'hFF;
            15'd12465: data <= 8'hFF;
            15'd12466: data <= 8'hFF;
            15'd12467: data <= 8'hFF;
            15'd12468: data <= 8'hFF;
            15'd12469: data <= 8'hF8;
            15'd12470: data <= 8'h0F;
            15'd12471: data <= 8'hFF;
            15'd12472: data <= 8'hFF;
            15'd12473: data <= 8'hFF;
            15'd12474: data <= 8'h80;
            15'd12475: data <= 8'h00;
            15'd12476: data <= 8'h00;
            15'd12477: data <= 8'h00;
            15'd12478: data <= 8'h00;
            15'd12479: data <= 8'h00;
            15'd12480: data <= 8'h00;
            15'd12481: data <= 8'h00;
            15'd12482: data <= 8'h00;
            15'd12483: data <= 8'h00;
            15'd12484: data <= 8'h00;
            15'd12485: data <= 8'h03;
            15'd12486: data <= 8'hFF;
            15'd12487: data <= 8'hFF;
            15'd12488: data <= 8'hC0;
            15'd12489: data <= 8'h7F;
            15'd12490: data <= 8'hFF;
            15'd12491: data <= 8'hFF;
            15'd12492: data <= 8'hFF;
            15'd12493: data <= 8'hFF;
            15'd12494: data <= 8'hFF;
            15'd12495: data <= 8'hFF;
            15'd12496: data <= 8'hFF;
            15'd12497: data <= 8'hFF;
            15'd12498: data <= 8'hFF;
            15'd12499: data <= 8'hF8;
            15'd12500: data <= 8'h0F;
            15'd12501: data <= 8'hFF;
            15'd12502: data <= 8'hFF;
            15'd12503: data <= 8'hFF;
            15'd12504: data <= 8'h80;
            15'd12505: data <= 8'h00;
            15'd12506: data <= 8'h00;
            15'd12507: data <= 8'h00;
            15'd12508: data <= 8'h00;
            15'd12509: data <= 8'h00;
            15'd12510: data <= 8'h00;
            15'd12511: data <= 8'h00;
            15'd12512: data <= 8'h00;
            15'd12513: data <= 8'h00;
            15'd12514: data <= 8'h00;
            15'd12515: data <= 8'h03;
            15'd12516: data <= 8'hFF;
            15'd12517: data <= 8'hFF;
            15'd12518: data <= 8'h80;
            15'd12519: data <= 8'h7F;
            15'd12520: data <= 8'hFF;
            15'd12521: data <= 8'hFF;
            15'd12522: data <= 8'hFF;
            15'd12523: data <= 8'hFF;
            15'd12524: data <= 8'hFF;
            15'd12525: data <= 8'hFF;
            15'd12526: data <= 8'hFF;
            15'd12527: data <= 8'hFF;
            15'd12528: data <= 8'hFF;
            15'd12529: data <= 8'hF8;
            15'd12530: data <= 8'h07;
            15'd12531: data <= 8'hFF;
            15'd12532: data <= 8'hFF;
            15'd12533: data <= 8'hFF;
            15'd12534: data <= 8'h80;
            15'd12535: data <= 8'h00;
            15'd12536: data <= 8'h00;
            15'd12537: data <= 8'h00;
            15'd12538: data <= 8'h00;
            15'd12539: data <= 8'h00;
            15'd12540: data <= 8'h00;
            15'd12541: data <= 8'h00;
            15'd12542: data <= 8'h00;
            15'd12543: data <= 8'h00;
            15'd12544: data <= 8'h00;
            15'd12545: data <= 8'h03;
            15'd12546: data <= 8'hFF;
            15'd12547: data <= 8'hFF;
            15'd12548: data <= 8'h80;
            15'd12549: data <= 8'hFF;
            15'd12550: data <= 8'hFF;
            15'd12551: data <= 8'hFF;
            15'd12552: data <= 8'hFF;
            15'd12553: data <= 8'hFF;
            15'd12554: data <= 8'hFF;
            15'd12555: data <= 8'hFF;
            15'd12556: data <= 8'hFF;
            15'd12557: data <= 8'hFF;
            15'd12558: data <= 8'hFF;
            15'd12559: data <= 8'hFC;
            15'd12560: data <= 8'h07;
            15'd12561: data <= 8'hFF;
            15'd12562: data <= 8'hFF;
            15'd12563: data <= 8'hFF;
            15'd12564: data <= 8'h80;
            15'd12565: data <= 8'h00;
            15'd12566: data <= 8'h00;
            15'd12567: data <= 8'h00;
            15'd12568: data <= 8'h00;
            15'd12569: data <= 8'h00;
            15'd12570: data <= 8'h00;
            15'd12571: data <= 8'h00;
            15'd12572: data <= 8'h00;
            15'd12573: data <= 8'h00;
            15'd12574: data <= 8'h00;
            15'd12575: data <= 8'h03;
            15'd12576: data <= 8'hFF;
            15'd12577: data <= 8'hFF;
            15'd12578: data <= 8'h00;
            15'd12579: data <= 8'hFF;
            15'd12580: data <= 8'hFF;
            15'd12581: data <= 8'hFF;
            15'd12582: data <= 8'hFF;
            15'd12583: data <= 8'hFF;
            15'd12584: data <= 8'hFF;
            15'd12585: data <= 8'hFF;
            15'd12586: data <= 8'hFF;
            15'd12587: data <= 8'hFF;
            15'd12588: data <= 8'hFF;
            15'd12589: data <= 8'hFC;
            15'd12590: data <= 8'h07;
            15'd12591: data <= 8'hFF;
            15'd12592: data <= 8'hFF;
            15'd12593: data <= 8'hFF;
            15'd12594: data <= 8'h80;
            15'd12595: data <= 8'h00;
            15'd12596: data <= 8'h00;
            15'd12597: data <= 8'h00;
            15'd12598: data <= 8'h00;
            15'd12599: data <= 8'h00;
            15'd12600: data <= 8'h00;
            15'd12601: data <= 8'h00;
            15'd12602: data <= 8'h00;
            15'd12603: data <= 8'h00;
            15'd12604: data <= 8'h00;
            15'd12605: data <= 8'h03;
            15'd12606: data <= 8'hFF;
            15'd12607: data <= 8'hFF;
            15'd12608: data <= 8'h01;
            15'd12609: data <= 8'hFF;
            15'd12610: data <= 8'hFF;
            15'd12611: data <= 8'hFF;
            15'd12612: data <= 8'hFF;
            15'd12613: data <= 8'hFF;
            15'd12614: data <= 8'hFF;
            15'd12615: data <= 8'hFF;
            15'd12616: data <= 8'hFF;
            15'd12617: data <= 8'hFF;
            15'd12618: data <= 8'hFF;
            15'd12619: data <= 8'hFE;
            15'd12620: data <= 8'h03;
            15'd12621: data <= 8'hFF;
            15'd12622: data <= 8'hFF;
            15'd12623: data <= 8'hFF;
            15'd12624: data <= 8'h80;
            15'd12625: data <= 8'h00;
            15'd12626: data <= 8'h00;
            15'd12627: data <= 8'h00;
            15'd12628: data <= 8'h00;
            15'd12629: data <= 8'h00;
            15'd12630: data <= 8'h00;
            15'd12631: data <= 8'h00;
            15'd12632: data <= 8'h00;
            15'd12633: data <= 8'h00;
            15'd12634: data <= 8'h00;
            15'd12635: data <= 8'h03;
            15'd12636: data <= 8'hFF;
            15'd12637: data <= 8'hFF;
            15'd12638: data <= 8'h01;
            15'd12639: data <= 8'hFF;
            15'd12640: data <= 8'hFF;
            15'd12641: data <= 8'hFF;
            15'd12642: data <= 8'hFF;
            15'd12643: data <= 8'hFF;
            15'd12644: data <= 8'hFF;
            15'd12645: data <= 8'hFF;
            15'd12646: data <= 8'hFF;
            15'd12647: data <= 8'hFF;
            15'd12648: data <= 8'hFF;
            15'd12649: data <= 8'hFE;
            15'd12650: data <= 8'h01;
            15'd12651: data <= 8'hFF;
            15'd12652: data <= 8'hFF;
            15'd12653: data <= 8'hFF;
            15'd12654: data <= 8'h80;
            15'd12655: data <= 8'h00;
            15'd12656: data <= 8'h00;
            15'd12657: data <= 8'h00;
            15'd12658: data <= 8'h00;
            15'd12659: data <= 8'h00;
            15'd12660: data <= 8'h00;
            15'd12661: data <= 8'h00;
            15'd12662: data <= 8'h00;
            15'd12663: data <= 8'h00;
            15'd12664: data <= 8'h00;
            15'd12665: data <= 8'h03;
            15'd12666: data <= 8'hFF;
            15'd12667: data <= 8'hFF;
            15'd12668: data <= 8'h01;
            15'd12669: data <= 8'hFF;
            15'd12670: data <= 8'hF9;
            15'd12671: data <= 8'hFF;
            15'd12672: data <= 8'hFF;
            15'd12673: data <= 8'hFF;
            15'd12674: data <= 8'hFF;
            15'd12675: data <= 8'hFF;
            15'd12676: data <= 8'hFF;
            15'd12677: data <= 8'hFF;
            15'd12678: data <= 8'hFF;
            15'd12679: data <= 8'hFE;
            15'd12680: data <= 8'h01;
            15'd12681: data <= 8'hFF;
            15'd12682: data <= 8'hFF;
            15'd12683: data <= 8'hFF;
            15'd12684: data <= 8'h80;
            15'd12685: data <= 8'h00;
            15'd12686: data <= 8'h00;
            15'd12687: data <= 8'h00;
            15'd12688: data <= 8'h00;
            15'd12689: data <= 8'h00;
            15'd12690: data <= 8'h00;
            15'd12691: data <= 8'h00;
            15'd12692: data <= 8'h00;
            15'd12693: data <= 8'h00;
            15'd12694: data <= 8'h00;
            15'd12695: data <= 8'h03;
            15'd12696: data <= 8'hFF;
            15'd12697: data <= 8'hFE;
            15'd12698: data <= 8'h03;
            15'd12699: data <= 8'hFF;
            15'd12700: data <= 8'hF0;
            15'd12701: data <= 8'hFF;
            15'd12702: data <= 8'hFF;
            15'd12703: data <= 8'hFF;
            15'd12704: data <= 8'hFF;
            15'd12705: data <= 8'hFF;
            15'd12706: data <= 8'hFF;
            15'd12707: data <= 8'hFF;
            15'd12708: data <= 8'hFF;
            15'd12709: data <= 8'hFF;
            15'd12710: data <= 8'h00;
            15'd12711: data <= 8'hFF;
            15'd12712: data <= 8'hFF;
            15'd12713: data <= 8'hFF;
            15'd12714: data <= 8'h80;
            15'd12715: data <= 8'h00;
            15'd12716: data <= 8'h00;
            15'd12717: data <= 8'h00;
            15'd12718: data <= 8'h00;
            15'd12719: data <= 8'h00;
            15'd12720: data <= 8'h00;
            15'd12721: data <= 8'h00;
            15'd12722: data <= 8'h00;
            15'd12723: data <= 8'h00;
            15'd12724: data <= 8'h00;
            15'd12725: data <= 8'h03;
            15'd12726: data <= 8'hFF;
            15'd12727: data <= 8'hFE;
            15'd12728: data <= 8'h03;
            15'd12729: data <= 8'hFF;
            15'd12730: data <= 8'hF0;
            15'd12731: data <= 8'hFF;
            15'd12732: data <= 8'hC7;
            15'd12733: data <= 8'hFF;
            15'd12734: data <= 8'hFF;
            15'd12735: data <= 8'hFF;
            15'd12736: data <= 8'hFF;
            15'd12737: data <= 8'hFF;
            15'd12738: data <= 8'hFF;
            15'd12739: data <= 8'hFF;
            15'd12740: data <= 8'h00;
            15'd12741: data <= 8'hFF;
            15'd12742: data <= 8'hFF;
            15'd12743: data <= 8'hFF;
            15'd12744: data <= 8'h80;
            15'd12745: data <= 8'h00;
            15'd12746: data <= 8'h00;
            15'd12747: data <= 8'h00;
            15'd12748: data <= 8'h00;
            15'd12749: data <= 8'h00;
            15'd12750: data <= 8'h00;
            15'd12751: data <= 8'h00;
            15'd12752: data <= 8'h00;
            15'd12753: data <= 8'h00;
            15'd12754: data <= 8'h00;
            15'd12755: data <= 8'h03;
            15'd12756: data <= 8'hFF;
            15'd12757: data <= 8'hFE;
            15'd12758: data <= 8'h07;
            15'd12759: data <= 8'hFF;
            15'd12760: data <= 8'hF0;
            15'd12761: data <= 8'hFF;
            15'd12762: data <= 8'h83;
            15'd12763: data <= 8'hFF;
            15'd12764: data <= 8'hFF;
            15'd12765: data <= 8'hFF;
            15'd12766: data <= 8'hFF;
            15'd12767: data <= 8'hFF;
            15'd12768: data <= 8'hFF;
            15'd12769: data <= 8'hFF;
            15'd12770: data <= 8'h80;
            15'd12771: data <= 8'h7F;
            15'd12772: data <= 8'hFF;
            15'd12773: data <= 8'hFF;
            15'd12774: data <= 8'h80;
            15'd12775: data <= 8'h00;
            15'd12776: data <= 8'h00;
            15'd12777: data <= 8'h00;
            15'd12778: data <= 8'h00;
            15'd12779: data <= 8'h00;
            15'd12780: data <= 8'h00;
            15'd12781: data <= 8'h00;
            15'd12782: data <= 8'h00;
            15'd12783: data <= 8'h00;
            15'd12784: data <= 8'h00;
            15'd12785: data <= 8'h03;
            15'd12786: data <= 8'hFF;
            15'd12787: data <= 8'hFE;
            15'd12788: data <= 8'h07;
            15'd12789: data <= 8'hFF;
            15'd12790: data <= 8'hFD;
            15'd12791: data <= 8'hFF;
            15'd12792: data <= 8'h83;
            15'd12793: data <= 8'hFF;
            15'd12794: data <= 8'hFF;
            15'd12795: data <= 8'hFF;
            15'd12796: data <= 8'hFF;
            15'd12797: data <= 8'hFF;
            15'd12798: data <= 8'hFF;
            15'd12799: data <= 8'hFF;
            15'd12800: data <= 8'h80;
            15'd12801: data <= 8'h7F;
            15'd12802: data <= 8'hFF;
            15'd12803: data <= 8'hFF;
            15'd12804: data <= 8'h80;
            15'd12805: data <= 8'h00;
            15'd12806: data <= 8'h00;
            15'd12807: data <= 8'h00;
            15'd12808: data <= 8'h00;
            15'd12809: data <= 8'h00;
            15'd12810: data <= 8'h00;
            15'd12811: data <= 8'h00;
            15'd12812: data <= 8'h00;
            15'd12813: data <= 8'h00;
            15'd12814: data <= 8'h00;
            15'd12815: data <= 8'h03;
            15'd12816: data <= 8'hFF;
            15'd12817: data <= 8'hFE;
            15'd12818: data <= 8'h07;
            15'd12819: data <= 8'hFF;
            15'd12820: data <= 8'hFF;
            15'd12821: data <= 8'hFF;
            15'd12822: data <= 8'h83;
            15'd12823: data <= 8'hFF;
            15'd12824: data <= 8'hFF;
            15'd12825: data <= 8'hFF;
            15'd12826: data <= 8'hFF;
            15'd12827: data <= 8'hFF;
            15'd12828: data <= 8'hFF;
            15'd12829: data <= 8'hFF;
            15'd12830: data <= 8'hC0;
            15'd12831: data <= 8'h3F;
            15'd12832: data <= 8'hFF;
            15'd12833: data <= 8'hFF;
            15'd12834: data <= 8'h80;
            15'd12835: data <= 8'h00;
            15'd12836: data <= 8'h00;
            15'd12837: data <= 8'h00;
            15'd12838: data <= 8'h00;
            15'd12839: data <= 8'h00;
            15'd12840: data <= 8'h00;
            15'd12841: data <= 8'h00;
            15'd12842: data <= 8'h00;
            15'd12843: data <= 8'h00;
            15'd12844: data <= 8'h00;
            15'd12845: data <= 8'h03;
            15'd12846: data <= 8'hFF;
            15'd12847: data <= 8'hFE;
            15'd12848: data <= 8'h07;
            15'd12849: data <= 8'hFF;
            15'd12850: data <= 8'hFF;
            15'd12851: data <= 8'hFF;
            15'd12852: data <= 8'hEF;
            15'd12853: data <= 8'hFF;
            15'd12854: data <= 8'hFF;
            15'd12855: data <= 8'hFF;
            15'd12856: data <= 8'hFF;
            15'd12857: data <= 8'hFF;
            15'd12858: data <= 8'hFF;
            15'd12859: data <= 8'hFF;
            15'd12860: data <= 8'hE0;
            15'd12861: data <= 8'h3F;
            15'd12862: data <= 8'hFF;
            15'd12863: data <= 8'hFF;
            15'd12864: data <= 8'h80;
            15'd12865: data <= 8'h00;
            15'd12866: data <= 8'h00;
            15'd12867: data <= 8'h00;
            15'd12868: data <= 8'h00;
            15'd12869: data <= 8'h00;
            15'd12870: data <= 8'h00;
            15'd12871: data <= 8'h00;
            15'd12872: data <= 8'h00;
            15'd12873: data <= 8'h00;
            15'd12874: data <= 8'h00;
            15'd12875: data <= 8'h03;
            15'd12876: data <= 8'hFF;
            15'd12877: data <= 8'hFE;
            15'd12878: data <= 8'h07;
            15'd12879: data <= 8'hFF;
            15'd12880: data <= 8'hFF;
            15'd12881: data <= 8'hFF;
            15'd12882: data <= 8'hFF;
            15'd12883: data <= 8'hFF;
            15'd12884: data <= 8'hFF;
            15'd12885: data <= 8'hFF;
            15'd12886: data <= 8'hFF;
            15'd12887: data <= 8'hFF;
            15'd12888: data <= 8'hFF;
            15'd12889: data <= 8'hFF;
            15'd12890: data <= 8'hE0;
            15'd12891: data <= 8'h1F;
            15'd12892: data <= 8'hFF;
            15'd12893: data <= 8'hFF;
            15'd12894: data <= 8'h80;
            15'd12895: data <= 8'h00;
            15'd12896: data <= 8'h00;
            15'd12897: data <= 8'h00;
            15'd12898: data <= 8'h00;
            15'd12899: data <= 8'h00;
            15'd12900: data <= 8'h00;
            15'd12901: data <= 8'h00;
            15'd12902: data <= 8'h00;
            15'd12903: data <= 8'h00;
            15'd12904: data <= 8'h00;
            15'd12905: data <= 8'h03;
            15'd12906: data <= 8'hFF;
            15'd12907: data <= 8'hFE;
            15'd12908: data <= 8'h07;
            15'd12909: data <= 8'hFF;
            15'd12910: data <= 8'hFF;
            15'd12911: data <= 8'hFF;
            15'd12912: data <= 8'hFF;
            15'd12913: data <= 8'hFF;
            15'd12914: data <= 8'hFF;
            15'd12915: data <= 8'hFF;
            15'd12916: data <= 8'hFF;
            15'd12917: data <= 8'hFF;
            15'd12918: data <= 8'hFF;
            15'd12919: data <= 8'hFF;
            15'd12920: data <= 8'hF0;
            15'd12921: data <= 8'h0F;
            15'd12922: data <= 8'hFF;
            15'd12923: data <= 8'hFF;
            15'd12924: data <= 8'h80;
            15'd12925: data <= 8'h00;
            15'd12926: data <= 8'h00;
            15'd12927: data <= 8'h00;
            15'd12928: data <= 8'h00;
            15'd12929: data <= 8'h00;
            15'd12930: data <= 8'h00;
            15'd12931: data <= 8'h00;
            15'd12932: data <= 8'h00;
            15'd12933: data <= 8'h00;
            15'd12934: data <= 8'h00;
            15'd12935: data <= 8'h03;
            15'd12936: data <= 8'hFF;
            15'd12937: data <= 8'hFE;
            15'd12938: data <= 8'h07;
            15'd12939: data <= 8'hFF;
            15'd12940: data <= 8'hFF;
            15'd12941: data <= 8'hFF;
            15'd12942: data <= 8'hFF;
            15'd12943: data <= 8'hFF;
            15'd12944: data <= 8'hFF;
            15'd12945: data <= 8'hFF;
            15'd12946: data <= 8'hFF;
            15'd12947: data <= 8'hFF;
            15'd12948: data <= 8'hFF;
            15'd12949: data <= 8'hFF;
            15'd12950: data <= 8'hF0;
            15'd12951: data <= 8'h0F;
            15'd12952: data <= 8'hFF;
            15'd12953: data <= 8'hFF;
            15'd12954: data <= 8'h80;
            15'd12955: data <= 8'h00;
            15'd12956: data <= 8'h00;
            15'd12957: data <= 8'h00;
            15'd12958: data <= 8'h00;
            15'd12959: data <= 8'h00;
            15'd12960: data <= 8'h00;
            15'd12961: data <= 8'h00;
            15'd12962: data <= 8'h00;
            15'd12963: data <= 8'h00;
            15'd12964: data <= 8'h00;
            15'd12965: data <= 8'h03;
            15'd12966: data <= 8'hFF;
            15'd12967: data <= 8'hFE;
            15'd12968: data <= 8'h07;
            15'd12969: data <= 8'hFF;
            15'd12970: data <= 8'hFF;
            15'd12971: data <= 8'hFF;
            15'd12972: data <= 8'hFF;
            15'd12973: data <= 8'hFF;
            15'd12974: data <= 8'hFF;
            15'd12975: data <= 8'hFF;
            15'd12976: data <= 8'hFF;
            15'd12977: data <= 8'hFF;
            15'd12978: data <= 8'hFF;
            15'd12979: data <= 8'hFF;
            15'd12980: data <= 8'hF8;
            15'd12981: data <= 8'h0F;
            15'd12982: data <= 8'hFF;
            15'd12983: data <= 8'hFF;
            15'd12984: data <= 8'h80;
            15'd12985: data <= 8'h00;
            15'd12986: data <= 8'h00;
            15'd12987: data <= 8'h00;
            15'd12988: data <= 8'h00;
            15'd12989: data <= 8'h00;
            15'd12990: data <= 8'h00;
            15'd12991: data <= 8'h00;
            15'd12992: data <= 8'h00;
            15'd12993: data <= 8'h00;
            15'd12994: data <= 8'h00;
            15'd12995: data <= 8'h03;
            15'd12996: data <= 8'hFF;
            15'd12997: data <= 8'hFE;
            15'd12998: data <= 8'h07;
            15'd12999: data <= 8'hFF;
            15'd13000: data <= 8'hFF;
            15'd13001: data <= 8'hFF;
            15'd13002: data <= 8'hFF;
            15'd13003: data <= 8'hFF;
            15'd13004: data <= 8'hFF;
            15'd13005: data <= 8'hFF;
            15'd13006: data <= 8'hFF;
            15'd13007: data <= 8'hFF;
            15'd13008: data <= 8'hFF;
            15'd13009: data <= 8'hFF;
            15'd13010: data <= 8'hFC;
            15'd13011: data <= 8'h07;
            15'd13012: data <= 8'hFF;
            15'd13013: data <= 8'hFF;
            15'd13014: data <= 8'h80;
            15'd13015: data <= 8'h00;
            15'd13016: data <= 8'h00;
            15'd13017: data <= 8'h00;
            15'd13018: data <= 8'h00;
            15'd13019: data <= 8'h00;
            15'd13020: data <= 8'h00;
            15'd13021: data <= 8'h00;
            15'd13022: data <= 8'h00;
            15'd13023: data <= 8'h00;
            15'd13024: data <= 8'h00;
            15'd13025: data <= 8'h03;
            15'd13026: data <= 8'hFF;
            15'd13027: data <= 8'hFE;
            15'd13028: data <= 8'h07;
            15'd13029: data <= 8'hFF;
            15'd13030: data <= 8'hFB;
            15'd13031: data <= 8'hFF;
            15'd13032: data <= 8'hFF;
            15'd13033: data <= 8'hFF;
            15'd13034: data <= 8'hFF;
            15'd13035: data <= 8'hFF;
            15'd13036: data <= 8'hFF;
            15'd13037: data <= 8'hFF;
            15'd13038: data <= 8'hFF;
            15'd13039: data <= 8'hFF;
            15'd13040: data <= 8'hFC;
            15'd13041: data <= 8'h07;
            15'd13042: data <= 8'hFF;
            15'd13043: data <= 8'hFF;
            15'd13044: data <= 8'h80;
            15'd13045: data <= 8'h00;
            15'd13046: data <= 8'h00;
            15'd13047: data <= 8'h00;
            15'd13048: data <= 8'h00;
            15'd13049: data <= 8'h00;
            15'd13050: data <= 8'h00;
            15'd13051: data <= 8'h00;
            15'd13052: data <= 8'h00;
            15'd13053: data <= 8'h00;
            15'd13054: data <= 8'h00;
            15'd13055: data <= 8'h03;
            15'd13056: data <= 8'hFF;
            15'd13057: data <= 8'hFF;
            15'd13058: data <= 8'h03;
            15'd13059: data <= 8'hFF;
            15'd13060: data <= 8'hF1;
            15'd13061: data <= 8'hFF;
            15'd13062: data <= 8'hFF;
            15'd13063: data <= 8'hFF;
            15'd13064: data <= 8'hFF;
            15'd13065: data <= 8'hFF;
            15'd13066: data <= 8'hFF;
            15'd13067: data <= 8'hFF;
            15'd13068: data <= 8'hFF;
            15'd13069: data <= 8'hFF;
            15'd13070: data <= 8'hFE;
            15'd13071: data <= 8'h03;
            15'd13072: data <= 8'hFF;
            15'd13073: data <= 8'hFF;
            15'd13074: data <= 8'h80;
            15'd13075: data <= 8'h00;
            15'd13076: data <= 8'h00;
            15'd13077: data <= 8'h00;
            15'd13078: data <= 8'h00;
            15'd13079: data <= 8'h00;
            15'd13080: data <= 8'h00;
            15'd13081: data <= 8'h00;
            15'd13082: data <= 8'h00;
            15'd13083: data <= 8'h00;
            15'd13084: data <= 8'h00;
            15'd13085: data <= 8'h03;
            15'd13086: data <= 8'hFF;
            15'd13087: data <= 8'hFF;
            15'd13088: data <= 8'h03;
            15'd13089: data <= 8'hFF;
            15'd13090: data <= 8'hE0;
            15'd13091: data <= 8'h38;
            15'd13092: data <= 8'h3F;
            15'd13093: data <= 8'hFF;
            15'd13094: data <= 8'hFF;
            15'd13095: data <= 8'hFF;
            15'd13096: data <= 8'hFF;
            15'd13097: data <= 8'hFF;
            15'd13098: data <= 8'hFF;
            15'd13099: data <= 8'hFF;
            15'd13100: data <= 8'hFE;
            15'd13101: data <= 8'h03;
            15'd13102: data <= 8'hFF;
            15'd13103: data <= 8'hFF;
            15'd13104: data <= 8'h80;
            15'd13105: data <= 8'h00;
            15'd13106: data <= 8'h00;
            15'd13107: data <= 8'h00;
            15'd13108: data <= 8'h00;
            15'd13109: data <= 8'h00;
            15'd13110: data <= 8'h00;
            15'd13111: data <= 8'h00;
            15'd13112: data <= 8'h00;
            15'd13113: data <= 8'h00;
            15'd13114: data <= 8'h00;
            15'd13115: data <= 8'h03;
            15'd13116: data <= 8'hFF;
            15'd13117: data <= 8'hFF;
            15'd13118: data <= 8'h83;
            15'd13119: data <= 8'hFF;
            15'd13120: data <= 8'hE0;
            15'd13121: data <= 8'h00;
            15'd13122: data <= 8'h3F;
            15'd13123: data <= 8'hFF;
            15'd13124: data <= 8'hFF;
            15'd13125: data <= 8'hFF;
            15'd13126: data <= 8'hFF;
            15'd13127: data <= 8'hFF;
            15'd13128: data <= 8'hFF;
            15'd13129: data <= 8'hFF;
            15'd13130: data <= 8'hFF;
            15'd13131: data <= 8'h01;
            15'd13132: data <= 8'hFF;
            15'd13133: data <= 8'hFF;
            15'd13134: data <= 8'h80;
            15'd13135: data <= 8'h00;
            15'd13136: data <= 8'h00;
            15'd13137: data <= 8'h00;
            15'd13138: data <= 8'h00;
            15'd13139: data <= 8'h00;
            15'd13140: data <= 8'h00;
            15'd13141: data <= 8'h00;
            15'd13142: data <= 8'h00;
            15'd13143: data <= 8'h00;
            15'd13144: data <= 8'h00;
            15'd13145: data <= 8'h03;
            15'd13146: data <= 8'hFF;
            15'd13147: data <= 8'hFF;
            15'd13148: data <= 8'h81;
            15'd13149: data <= 8'h03;
            15'd13150: data <= 8'hE0;
            15'd13151: data <= 8'h00;
            15'd13152: data <= 8'h3F;
            15'd13153: data <= 8'hFF;
            15'd13154: data <= 8'hFF;
            15'd13155: data <= 8'hFF;
            15'd13156: data <= 8'hFF;
            15'd13157: data <= 8'hFF;
            15'd13158: data <= 8'hFF;
            15'd13159: data <= 8'hFF;
            15'd13160: data <= 8'hFF;
            15'd13161: data <= 8'h00;
            15'd13162: data <= 8'hFF;
            15'd13163: data <= 8'hFF;
            15'd13164: data <= 8'h80;
            15'd13165: data <= 8'h00;
            15'd13166: data <= 8'h00;
            15'd13167: data <= 8'h00;
            15'd13168: data <= 8'h00;
            15'd13169: data <= 8'h00;
            15'd13170: data <= 8'h00;
            15'd13171: data <= 8'h00;
            15'd13172: data <= 8'h00;
            15'd13173: data <= 8'h00;
            15'd13174: data <= 8'h00;
            15'd13175: data <= 8'h03;
            15'd13176: data <= 8'hFF;
            15'd13177: data <= 8'hFF;
            15'd13178: data <= 8'hC0;
            15'd13179: data <= 8'h00;
            15'd13180: data <= 8'h70;
            15'd13181: data <= 8'h00;
            15'd13182: data <= 8'h1F;
            15'd13183: data <= 8'hFF;
            15'd13184: data <= 8'hFF;
            15'd13185: data <= 8'hFF;
            15'd13186: data <= 8'hFF;
            15'd13187: data <= 8'hFF;
            15'd13188: data <= 8'hFF;
            15'd13189: data <= 8'hFF;
            15'd13190: data <= 8'hFF;
            15'd13191: data <= 8'h80;
            15'd13192: data <= 8'h7F;
            15'd13193: data <= 8'hFF;
            15'd13194: data <= 8'h80;
            15'd13195: data <= 8'h00;
            15'd13196: data <= 8'h00;
            15'd13197: data <= 8'h00;
            15'd13198: data <= 8'h00;
            15'd13199: data <= 8'h00;
            15'd13200: data <= 8'h00;
            15'd13201: data <= 8'h00;
            15'd13202: data <= 8'h00;
            15'd13203: data <= 8'h00;
            15'd13204: data <= 8'h00;
            15'd13205: data <= 8'h03;
            15'd13206: data <= 8'hFF;
            15'd13207: data <= 8'hFF;
            15'd13208: data <= 8'hE0;
            15'd13209: data <= 8'h00;
            15'd13210: data <= 8'h18;
            15'd13211: data <= 8'h00;
            15'd13212: data <= 8'h7F;
            15'd13213: data <= 8'hFF;
            15'd13214: data <= 8'hFF;
            15'd13215: data <= 8'hFF;
            15'd13216: data <= 8'hFF;
            15'd13217: data <= 8'hFF;
            15'd13218: data <= 8'hFF;
            15'd13219: data <= 8'hFF;
            15'd13220: data <= 8'hFF;
            15'd13221: data <= 8'h80;
            15'd13222: data <= 8'h7F;
            15'd13223: data <= 8'hFF;
            15'd13224: data <= 8'h80;
            15'd13225: data <= 8'h00;
            15'd13226: data <= 8'h00;
            15'd13227: data <= 8'h00;
            15'd13228: data <= 8'h00;
            15'd13229: data <= 8'h00;
            15'd13230: data <= 8'h00;
            15'd13231: data <= 8'h00;
            15'd13232: data <= 8'h00;
            15'd13233: data <= 8'h00;
            15'd13234: data <= 8'h00;
            15'd13235: data <= 8'h03;
            15'd13236: data <= 8'hFF;
            15'd13237: data <= 8'hFF;
            15'd13238: data <= 8'hC0;
            15'd13239: data <= 8'h00;
            15'd13240: data <= 8'h03;
            15'd13241: data <= 8'hF3;
            15'd13242: data <= 8'hFF;
            15'd13243: data <= 8'hFF;
            15'd13244: data <= 8'hFF;
            15'd13245: data <= 8'hFF;
            15'd13246: data <= 8'hFF;
            15'd13247: data <= 8'hFF;
            15'd13248: data <= 8'hFF;
            15'd13249: data <= 8'hFF;
            15'd13250: data <= 8'hFF;
            15'd13251: data <= 8'hC0;
            15'd13252: data <= 8'h7F;
            15'd13253: data <= 8'hFF;
            15'd13254: data <= 8'h80;
            15'd13255: data <= 8'h00;
            15'd13256: data <= 8'h00;
            15'd13257: data <= 8'h00;
            15'd13258: data <= 8'h00;
            15'd13259: data <= 8'h00;
            15'd13260: data <= 8'h00;
            15'd13261: data <= 8'h00;
            15'd13262: data <= 8'h00;
            15'd13263: data <= 8'h00;
            15'd13264: data <= 8'h00;
            15'd13265: data <= 8'h03;
            15'd13266: data <= 8'hFF;
            15'd13267: data <= 8'hFF;
            15'd13268: data <= 8'hC0;
            15'd13269: data <= 8'h00;
            15'd13270: data <= 8'h01;
            15'd13271: data <= 8'hFF;
            15'd13272: data <= 8'hF8;
            15'd13273: data <= 8'h7F;
            15'd13274: data <= 8'hFF;
            15'd13275: data <= 8'hFF;
            15'd13276: data <= 8'hFF;
            15'd13277: data <= 8'hFF;
            15'd13278: data <= 8'hFF;
            15'd13279: data <= 8'hFF;
            15'd13280: data <= 8'hFF;
            15'd13281: data <= 8'hC0;
            15'd13282: data <= 8'h3F;
            15'd13283: data <= 8'hFF;
            15'd13284: data <= 8'h80;
            15'd13285: data <= 8'h00;
            15'd13286: data <= 8'h00;
            15'd13287: data <= 8'h00;
            15'd13288: data <= 8'h00;
            15'd13289: data <= 8'h00;
            15'd13290: data <= 8'h00;
            15'd13291: data <= 8'h00;
            15'd13292: data <= 8'h00;
            15'd13293: data <= 8'h00;
            15'd13294: data <= 8'h00;
            15'd13295: data <= 8'h03;
            15'd13296: data <= 8'hFF;
            15'd13297: data <= 8'hFF;
            15'd13298: data <= 8'hF0;
            15'd13299: data <= 8'h00;
            15'd13300: data <= 8'h00;
            15'd13301: data <= 8'h0F;
            15'd13302: data <= 8'hC0;
            15'd13303: data <= 8'h7F;
            15'd13304: data <= 8'hFF;
            15'd13305: data <= 8'hFF;
            15'd13306: data <= 8'hFF;
            15'd13307: data <= 8'hFF;
            15'd13308: data <= 8'hFF;
            15'd13309: data <= 8'hFF;
            15'd13310: data <= 8'hFF;
            15'd13311: data <= 8'hE0;
            15'd13312: data <= 8'h3F;
            15'd13313: data <= 8'hFF;
            15'd13314: data <= 8'h80;
            15'd13315: data <= 8'h00;
            15'd13316: data <= 8'h00;
            15'd13317: data <= 8'h00;
            15'd13318: data <= 8'h00;
            15'd13319: data <= 8'h00;
            15'd13320: data <= 8'h00;
            15'd13321: data <= 8'h00;
            15'd13322: data <= 8'h00;
            15'd13323: data <= 8'h00;
            15'd13324: data <= 8'h00;
            15'd13325: data <= 8'h03;
            15'd13326: data <= 8'hFF;
            15'd13327: data <= 8'hFF;
            15'd13328: data <= 8'hF8;
            15'd13329: data <= 8'h00;
            15'd13330: data <= 8'h00;
            15'd13331: data <= 8'h04;
            15'd13332: data <= 8'h00;
            15'd13333: data <= 8'h7F;
            15'd13334: data <= 8'hFF;
            15'd13335: data <= 8'hFF;
            15'd13336: data <= 8'hFF;
            15'd13337: data <= 8'hFF;
            15'd13338: data <= 8'hFF;
            15'd13339: data <= 8'hFF;
            15'd13340: data <= 8'hFF;
            15'd13341: data <= 8'hE0;
            15'd13342: data <= 8'h1F;
            15'd13343: data <= 8'hFF;
            15'd13344: data <= 8'h80;
            15'd13345: data <= 8'h00;
            15'd13346: data <= 8'h00;
            15'd13347: data <= 8'h00;
            15'd13348: data <= 8'h00;
            15'd13349: data <= 8'h00;
            15'd13350: data <= 8'h00;
            15'd13351: data <= 8'h00;
            15'd13352: data <= 8'h00;
            15'd13353: data <= 8'h00;
            15'd13354: data <= 8'h00;
            15'd13355: data <= 8'h03;
            15'd13356: data <= 8'hFF;
            15'd13357: data <= 8'hFF;
            15'd13358: data <= 8'hF8;
            15'd13359: data <= 8'h00;
            15'd13360: data <= 8'h00;
            15'd13361: data <= 8'h00;
            15'd13362: data <= 8'h00;
            15'd13363: data <= 8'hFF;
            15'd13364: data <= 8'hFF;
            15'd13365: data <= 8'hFF;
            15'd13366: data <= 8'hFF;
            15'd13367: data <= 8'hFF;
            15'd13368: data <= 8'hFF;
            15'd13369: data <= 8'hFF;
            15'd13370: data <= 8'hFF;
            15'd13371: data <= 8'hF0;
            15'd13372: data <= 8'h1F;
            15'd13373: data <= 8'hFF;
            15'd13374: data <= 8'h80;
            15'd13375: data <= 8'h00;
            15'd13376: data <= 8'h00;
            15'd13377: data <= 8'h00;
            15'd13378: data <= 8'h00;
            15'd13379: data <= 8'h00;
            15'd13380: data <= 8'h00;
            15'd13381: data <= 8'h00;
            15'd13382: data <= 8'h00;
            15'd13383: data <= 8'h00;
            15'd13384: data <= 8'h00;
            15'd13385: data <= 8'h03;
            15'd13386: data <= 8'hFF;
            15'd13387: data <= 8'hFF;
            15'd13388: data <= 8'hFE;
            15'd13389: data <= 8'h00;
            15'd13390: data <= 8'h08;
            15'd13391: data <= 8'h00;
            15'd13392: data <= 8'h01;
            15'd13393: data <= 8'hFF;
            15'd13394: data <= 8'hFF;
            15'd13395: data <= 8'hFF;
            15'd13396: data <= 8'hFF;
            15'd13397: data <= 8'hFF;
            15'd13398: data <= 8'hFF;
            15'd13399: data <= 8'hFF;
            15'd13400: data <= 8'hFF;
            15'd13401: data <= 8'hF0;
            15'd13402: data <= 8'h1F;
            15'd13403: data <= 8'hFF;
            15'd13404: data <= 8'h80;
            15'd13405: data <= 8'h00;
            15'd13406: data <= 8'h00;
            15'd13407: data <= 8'h00;
            15'd13408: data <= 8'h00;
            15'd13409: data <= 8'h00;
            15'd13410: data <= 8'h00;
            15'd13411: data <= 8'h00;
            15'd13412: data <= 8'h00;
            15'd13413: data <= 8'h00;
            15'd13414: data <= 8'h00;
            15'd13415: data <= 8'h03;
            15'd13416: data <= 8'hFF;
            15'd13417: data <= 8'hFF;
            15'd13418: data <= 8'hFF;
            15'd13419: data <= 8'h00;
            15'd13420: data <= 8'h04;
            15'd13421: data <= 8'h00;
            15'd13422: data <= 8'h01;
            15'd13423: data <= 8'hFF;
            15'd13424: data <= 8'hFF;
            15'd13425: data <= 8'hFF;
            15'd13426: data <= 8'hFF;
            15'd13427: data <= 8'hFF;
            15'd13428: data <= 8'hFF;
            15'd13429: data <= 8'hFF;
            15'd13430: data <= 8'hFF;
            15'd13431: data <= 8'hF8;
            15'd13432: data <= 8'h0F;
            15'd13433: data <= 8'hFF;
            15'd13434: data <= 8'h80;
            15'd13435: data <= 8'h00;
            15'd13436: data <= 8'h00;
            15'd13437: data <= 8'h00;
            15'd13438: data <= 8'h00;
            15'd13439: data <= 8'h00;
            15'd13440: data <= 8'h00;
            15'd13441: data <= 8'h00;
            15'd13442: data <= 8'h00;
            15'd13443: data <= 8'h00;
            15'd13444: data <= 8'h00;
            15'd13445: data <= 8'h03;
            15'd13446: data <= 8'hFF;
            15'd13447: data <= 8'hFF;
            15'd13448: data <= 8'hFF;
            15'd13449: data <= 8'h80;
            15'd13450: data <= 8'h07;
            15'd13451: data <= 8'h80;
            15'd13452: data <= 8'h03;
            15'd13453: data <= 8'hFF;
            15'd13454: data <= 8'hFF;
            15'd13455: data <= 8'hFF;
            15'd13456: data <= 8'hFF;
            15'd13457: data <= 8'hFF;
            15'd13458: data <= 8'hFF;
            15'd13459: data <= 8'hFF;
            15'd13460: data <= 8'hFF;
            15'd13461: data <= 8'hF8;
            15'd13462: data <= 8'h0F;
            15'd13463: data <= 8'hFF;
            15'd13464: data <= 8'h80;
            15'd13465: data <= 8'h00;
            15'd13466: data <= 8'h00;
            15'd13467: data <= 8'h00;
            15'd13468: data <= 8'h00;
            15'd13469: data <= 8'h00;
            15'd13470: data <= 8'h00;
            15'd13471: data <= 8'h00;
            15'd13472: data <= 8'h00;
            15'd13473: data <= 8'h00;
            15'd13474: data <= 8'h00;
            15'd13475: data <= 8'h03;
            15'd13476: data <= 8'hFF;
            15'd13477: data <= 8'hFF;
            15'd13478: data <= 8'hFF;
            15'd13479: data <= 8'hE0;
            15'd13480: data <= 8'h07;
            15'd13481: data <= 8'hFF;
            15'd13482: data <= 8'hC7;
            15'd13483: data <= 8'hFF;
            15'd13484: data <= 8'hFF;
            15'd13485: data <= 8'hFF;
            15'd13486: data <= 8'hFF;
            15'd13487: data <= 8'hFF;
            15'd13488: data <= 8'hFF;
            15'd13489: data <= 8'hFF;
            15'd13490: data <= 8'hFF;
            15'd13491: data <= 8'hFC;
            15'd13492: data <= 8'h07;
            15'd13493: data <= 8'hFF;
            15'd13494: data <= 8'h80;
            15'd13495: data <= 8'h00;
            15'd13496: data <= 8'h00;
            15'd13497: data <= 8'h00;
            15'd13498: data <= 8'h00;
            15'd13499: data <= 8'h00;
            15'd13500: data <= 8'h00;
            15'd13501: data <= 8'h00;
            15'd13502: data <= 8'h00;
            15'd13503: data <= 8'h00;
            15'd13504: data <= 8'h00;
            15'd13505: data <= 8'h03;
            15'd13506: data <= 8'hFF;
            15'd13507: data <= 8'hFF;
            15'd13508: data <= 8'hFF;
            15'd13509: data <= 8'hF0;
            15'd13510: data <= 8'h83;
            15'd13511: data <= 8'hFF;
            15'd13512: data <= 8'hC7;
            15'd13513: data <= 8'hFF;
            15'd13514: data <= 8'hFF;
            15'd13515: data <= 8'hFF;
            15'd13516: data <= 8'hFF;
            15'd13517: data <= 8'hFF;
            15'd13518: data <= 8'hFF;
            15'd13519: data <= 8'hFF;
            15'd13520: data <= 8'hFF;
            15'd13521: data <= 8'hFC;
            15'd13522: data <= 8'h07;
            15'd13523: data <= 8'hFF;
            15'd13524: data <= 8'h80;
            15'd13525: data <= 8'h00;
            15'd13526: data <= 8'h00;
            15'd13527: data <= 8'h00;
            15'd13528: data <= 8'h00;
            15'd13529: data <= 8'h00;
            15'd13530: data <= 8'h00;
            15'd13531: data <= 8'h00;
            15'd13532: data <= 8'h00;
            15'd13533: data <= 8'h00;
            15'd13534: data <= 8'h00;
            15'd13535: data <= 8'h03;
            15'd13536: data <= 8'hFF;
            15'd13537: data <= 8'hFF;
            15'd13538: data <= 8'hFF;
            15'd13539: data <= 8'hF0;
            15'd13540: data <= 8'hC1;
            15'd13541: data <= 8'hFF;
            15'd13542: data <= 8'hC7;
            15'd13543: data <= 8'hFF;
            15'd13544: data <= 8'hFF;
            15'd13545: data <= 8'hFF;
            15'd13546: data <= 8'hFF;
            15'd13547: data <= 8'hFF;
            15'd13548: data <= 8'hFF;
            15'd13549: data <= 8'hFF;
            15'd13550: data <= 8'hFF;
            15'd13551: data <= 8'hFC;
            15'd13552: data <= 8'h07;
            15'd13553: data <= 8'hFF;
            15'd13554: data <= 8'h80;
            15'd13555: data <= 8'h00;
            15'd13556: data <= 8'h00;
            15'd13557: data <= 8'h00;
            15'd13558: data <= 8'h00;
            15'd13559: data <= 8'h00;
            15'd13560: data <= 8'h00;
            15'd13561: data <= 8'h00;
            15'd13562: data <= 8'h00;
            15'd13563: data <= 8'h00;
            15'd13564: data <= 8'h00;
            15'd13565: data <= 8'h03;
            15'd13566: data <= 8'hFF;
            15'd13567: data <= 8'hFF;
            15'd13568: data <= 8'hFF;
            15'd13569: data <= 8'hF0;
            15'd13570: data <= 8'hE1;
            15'd13571: data <= 8'hFF;
            15'd13572: data <= 8'hC7;
            15'd13573: data <= 8'hFF;
            15'd13574: data <= 8'hFF;
            15'd13575: data <= 8'hFF;
            15'd13576: data <= 8'hFF;
            15'd13577: data <= 8'hFF;
            15'd13578: data <= 8'hFF;
            15'd13579: data <= 8'hFF;
            15'd13580: data <= 8'hFF;
            15'd13581: data <= 8'hFE;
            15'd13582: data <= 8'h03;
            15'd13583: data <= 8'hFF;
            15'd13584: data <= 8'h80;
            15'd13585: data <= 8'h00;
            15'd13586: data <= 8'h00;
            15'd13587: data <= 8'h00;
            15'd13588: data <= 8'h00;
            15'd13589: data <= 8'h00;
            15'd13590: data <= 8'h00;
            15'd13591: data <= 8'h00;
            15'd13592: data <= 8'h00;
            15'd13593: data <= 8'h00;
            15'd13594: data <= 8'h00;
            15'd13595: data <= 8'h03;
            15'd13596: data <= 8'hFF;
            15'd13597: data <= 8'hFF;
            15'd13598: data <= 8'hFF;
            15'd13599: data <= 8'hF0;
            15'd13600: data <= 8'hF0;
            15'd13601: data <= 8'hFF;
            15'd13602: data <= 8'hC7;
            15'd13603: data <= 8'hFF;
            15'd13604: data <= 8'hFF;
            15'd13605: data <= 8'hFF;
            15'd13606: data <= 8'hFF;
            15'd13607: data <= 8'hFF;
            15'd13608: data <= 8'hFF;
            15'd13609: data <= 8'hFF;
            15'd13610: data <= 8'hFF;
            15'd13611: data <= 8'hFE;
            15'd13612: data <= 8'h03;
            15'd13613: data <= 8'hFF;
            15'd13614: data <= 8'h80;
            15'd13615: data <= 8'h00;
            15'd13616: data <= 8'h00;
            15'd13617: data <= 8'h00;
            15'd13618: data <= 8'h00;
            15'd13619: data <= 8'h00;
            15'd13620: data <= 8'h00;
            15'd13621: data <= 8'h00;
            15'd13622: data <= 8'h00;
            15'd13623: data <= 8'h00;
            15'd13624: data <= 8'h00;
            15'd13625: data <= 8'h03;
            15'd13626: data <= 8'hFF;
            15'd13627: data <= 8'hFF;
            15'd13628: data <= 8'hFF;
            15'd13629: data <= 8'hF8;
            15'd13630: data <= 8'h70;
            15'd13631: data <= 8'hFF;
            15'd13632: data <= 8'hE3;
            15'd13633: data <= 8'hFF;
            15'd13634: data <= 8'hFF;
            15'd13635: data <= 8'hFF;
            15'd13636: data <= 8'hFF;
            15'd13637: data <= 8'hFF;
            15'd13638: data <= 8'hFF;
            15'd13639: data <= 8'hFF;
            15'd13640: data <= 8'hFF;
            15'd13641: data <= 8'hFF;
            15'd13642: data <= 8'h01;
            15'd13643: data <= 8'hFF;
            15'd13644: data <= 8'h80;
            15'd13645: data <= 8'h00;
            15'd13646: data <= 8'h00;
            15'd13647: data <= 8'h00;
            15'd13648: data <= 8'h00;
            15'd13649: data <= 8'h00;
            15'd13650: data <= 8'h00;
            15'd13651: data <= 8'h00;
            15'd13652: data <= 8'h00;
            15'd13653: data <= 8'h00;
            15'd13654: data <= 8'h00;
            15'd13655: data <= 8'h03;
            15'd13656: data <= 8'hFF;
            15'd13657: data <= 8'hFF;
            15'd13658: data <= 8'hFF;
            15'd13659: data <= 8'hF0;
            15'd13660: data <= 8'h78;
            15'd13661: data <= 8'hFF;
            15'd13662: data <= 8'hE1;
            15'd13663: data <= 8'hFF;
            15'd13664: data <= 8'hFF;
            15'd13665: data <= 8'hFF;
            15'd13666: data <= 8'hFF;
            15'd13667: data <= 8'hFF;
            15'd13668: data <= 8'hFF;
            15'd13669: data <= 8'hFF;
            15'd13670: data <= 8'hFF;
            15'd13671: data <= 8'hFF;
            15'd13672: data <= 8'h01;
            15'd13673: data <= 8'hFF;
            15'd13674: data <= 8'h80;
            15'd13675: data <= 8'h00;
            15'd13676: data <= 8'h00;
            15'd13677: data <= 8'h00;
            15'd13678: data <= 8'h00;
            15'd13679: data <= 8'h00;
            15'd13680: data <= 8'h00;
            15'd13681: data <= 8'h00;
            15'd13682: data <= 8'h00;
            15'd13683: data <= 8'h00;
            15'd13684: data <= 8'h00;
            15'd13685: data <= 8'h03;
            15'd13686: data <= 8'hFF;
            15'd13687: data <= 8'hFF;
            15'd13688: data <= 8'hFF;
            15'd13689: data <= 8'hF0;
            15'd13690: data <= 8'h78;
            15'd13691: data <= 8'h7F;
            15'd13692: data <= 8'hE0;
            15'd13693: data <= 8'hFF;
            15'd13694: data <= 8'hFF;
            15'd13695: data <= 8'hFF;
            15'd13696: data <= 8'hFF;
            15'd13697: data <= 8'hFF;
            15'd13698: data <= 8'hFF;
            15'd13699: data <= 8'hFF;
            15'd13700: data <= 8'hFF;
            15'd13701: data <= 8'hFF;
            15'd13702: data <= 8'h80;
            15'd13703: data <= 8'hFF;
            15'd13704: data <= 8'h80;
            15'd13705: data <= 8'h00;
            15'd13706: data <= 8'h00;
            15'd13707: data <= 8'h00;
            15'd13708: data <= 8'h00;
            15'd13709: data <= 8'h00;
            15'd13710: data <= 8'h00;
            15'd13711: data <= 8'h00;
            15'd13712: data <= 8'h00;
            15'd13713: data <= 8'h00;
            15'd13714: data <= 8'h00;
            15'd13715: data <= 8'h03;
            15'd13716: data <= 8'hFF;
            15'd13717: data <= 8'hFF;
            15'd13718: data <= 8'hFF;
            15'd13719: data <= 8'hF0;
            15'd13720: data <= 8'h78;
            15'd13721: data <= 8'h7F;
            15'd13722: data <= 8'hE0;
            15'd13723: data <= 8'h7F;
            15'd13724: data <= 8'hFF;
            15'd13725: data <= 8'hFF;
            15'd13726: data <= 8'hFF;
            15'd13727: data <= 8'hFF;
            15'd13728: data <= 8'hFF;
            15'd13729: data <= 8'hFF;
            15'd13730: data <= 8'hFF;
            15'd13731: data <= 8'hFF;
            15'd13732: data <= 8'h80;
            15'd13733: data <= 8'hFF;
            15'd13734: data <= 8'h80;
            15'd13735: data <= 8'h00;
            15'd13736: data <= 8'h00;
            15'd13737: data <= 8'h00;
            15'd13738: data <= 8'h00;
            15'd13739: data <= 8'h00;
            15'd13740: data <= 8'h00;
            15'd13741: data <= 8'h00;
            15'd13742: data <= 8'h00;
            15'd13743: data <= 8'h00;
            15'd13744: data <= 8'h00;
            15'd13745: data <= 8'h03;
            15'd13746: data <= 8'hFF;
            15'd13747: data <= 8'hFF;
            15'd13748: data <= 8'hFF;
            15'd13749: data <= 8'hF0;
            15'd13750: data <= 8'h7C;
            15'd13751: data <= 8'h3F;
            15'd13752: data <= 8'hF0;
            15'd13753: data <= 8'h3F;
            15'd13754: data <= 8'hFF;
            15'd13755: data <= 8'hFF;
            15'd13756: data <= 8'hF0;
            15'd13757: data <= 8'h7F;
            15'd13758: data <= 8'hFF;
            15'd13759: data <= 8'hFF;
            15'd13760: data <= 8'hFF;
            15'd13761: data <= 8'hFF;
            15'd13762: data <= 8'hC0;
            15'd13763: data <= 8'h7F;
            15'd13764: data <= 8'h80;
            15'd13765: data <= 8'h00;
            15'd13766: data <= 8'h00;
            15'd13767: data <= 8'h00;
            15'd13768: data <= 8'h00;
            15'd13769: data <= 8'h00;
            15'd13770: data <= 8'h00;
            15'd13771: data <= 8'h00;
            15'd13772: data <= 8'h00;
            15'd13773: data <= 8'h00;
            15'd13774: data <= 8'h00;
            15'd13775: data <= 8'h03;
            15'd13776: data <= 8'hFF;
            15'd13777: data <= 8'hFF;
            15'd13778: data <= 8'hFF;
            15'd13779: data <= 8'hF8;
            15'd13780: data <= 8'h7C;
            15'd13781: data <= 8'h3F;
            15'd13782: data <= 8'hF8;
            15'd13783: data <= 8'h0F;
            15'd13784: data <= 8'hFF;
            15'd13785: data <= 8'hFF;
            15'd13786: data <= 8'hE0;
            15'd13787: data <= 8'h7F;
            15'd13788: data <= 8'hFF;
            15'd13789: data <= 8'hFF;
            15'd13790: data <= 8'hFF;
            15'd13791: data <= 8'hFF;
            15'd13792: data <= 8'hC0;
            15'd13793: data <= 8'h7F;
            15'd13794: data <= 8'h80;
            15'd13795: data <= 8'h00;
            15'd13796: data <= 8'h00;
            15'd13797: data <= 8'h00;
            15'd13798: data <= 8'h00;
            15'd13799: data <= 8'h00;
            15'd13800: data <= 8'h00;
            15'd13801: data <= 8'h00;
            15'd13802: data <= 8'h00;
            15'd13803: data <= 8'h00;
            15'd13804: data <= 8'h00;
            15'd13805: data <= 8'h03;
            15'd13806: data <= 8'hFF;
            15'd13807: data <= 8'hFF;
            15'd13808: data <= 8'hFF;
            15'd13809: data <= 8'hF8;
            15'd13810: data <= 8'h7C;
            15'd13811: data <= 8'h3F;
            15'd13812: data <= 8'hFC;
            15'd13813: data <= 8'h03;
            15'd13814: data <= 8'hFF;
            15'd13815: data <= 8'hFF;
            15'd13816: data <= 8'hC0;
            15'd13817: data <= 8'h7F;
            15'd13818: data <= 8'hFF;
            15'd13819: data <= 8'hFF;
            15'd13820: data <= 8'hFF;
            15'd13821: data <= 8'hFF;
            15'd13822: data <= 8'hC0;
            15'd13823: data <= 8'h7F;
            15'd13824: data <= 8'h80;
            15'd13825: data <= 8'h00;
            15'd13826: data <= 8'h00;
            15'd13827: data <= 8'h00;
            15'd13828: data <= 8'h00;
            15'd13829: data <= 8'h00;
            15'd13830: data <= 8'h00;
            15'd13831: data <= 8'h00;
            15'd13832: data <= 8'h00;
            15'd13833: data <= 8'h00;
            15'd13834: data <= 8'h00;
            15'd13835: data <= 8'h03;
            15'd13836: data <= 8'hFF;
            15'd13837: data <= 8'hFF;
            15'd13838: data <= 8'hFF;
            15'd13839: data <= 8'hFC;
            15'd13840: data <= 8'h7C;
            15'd13841: data <= 8'h3F;
            15'd13842: data <= 8'hFE;
            15'd13843: data <= 8'h00;
            15'd13844: data <= 8'hFF;
            15'd13845: data <= 8'hFF;
            15'd13846: data <= 8'h00;
            15'd13847: data <= 8'h7F;
            15'd13848: data <= 8'hFF;
            15'd13849: data <= 8'hFF;
            15'd13850: data <= 8'hFF;
            15'd13851: data <= 8'hFF;
            15'd13852: data <= 8'hE0;
            15'd13853: data <= 8'h3F;
            15'd13854: data <= 8'h80;
            15'd13855: data <= 8'h00;
            15'd13856: data <= 8'h00;
            15'd13857: data <= 8'h00;
            15'd13858: data <= 8'h00;
            15'd13859: data <= 8'h00;
            15'd13860: data <= 8'h00;
            15'd13861: data <= 8'h00;
            15'd13862: data <= 8'h00;
            15'd13863: data <= 8'h00;
            15'd13864: data <= 8'h00;
            15'd13865: data <= 8'h03;
            15'd13866: data <= 8'hFF;
            15'd13867: data <= 8'hFF;
            15'd13868: data <= 8'hFF;
            15'd13869: data <= 8'hFC;
            15'd13870: data <= 8'h7C;
            15'd13871: data <= 8'h1F;
            15'd13872: data <= 8'hFF;
            15'd13873: data <= 8'h80;
            15'd13874: data <= 8'h1F;
            15'd13875: data <= 8'hFE;
            15'd13876: data <= 8'h00;
            15'd13877: data <= 8'h7F;
            15'd13878: data <= 8'hFF;
            15'd13879: data <= 8'hFF;
            15'd13880: data <= 8'hFF;
            15'd13881: data <= 8'hFF;
            15'd13882: data <= 8'hE0;
            15'd13883: data <= 8'h3F;
            15'd13884: data <= 8'h80;
            15'd13885: data <= 8'h00;
            15'd13886: data <= 8'h00;
            15'd13887: data <= 8'h00;
            15'd13888: data <= 8'h00;
            15'd13889: data <= 8'h00;
            15'd13890: data <= 8'h00;
            15'd13891: data <= 8'h00;
            15'd13892: data <= 8'h00;
            15'd13893: data <= 8'h00;
            15'd13894: data <= 8'h00;
            15'd13895: data <= 8'h03;
            15'd13896: data <= 8'hFF;
            15'd13897: data <= 8'hFF;
            15'd13898: data <= 8'hFF;
            15'd13899: data <= 8'hF8;
            15'd13900: data <= 8'h7E;
            15'd13901: data <= 8'h1F;
            15'd13902: data <= 8'hFF;
            15'd13903: data <= 8'hC0;
            15'd13904: data <= 8'h03;
            15'd13905: data <= 8'h00;
            15'd13906: data <= 8'h00;
            15'd13907: data <= 8'hFF;
            15'd13908: data <= 8'hFF;
            15'd13909: data <= 8'hFF;
            15'd13910: data <= 8'hFF;
            15'd13911: data <= 8'hFF;
            15'd13912: data <= 8'hE0;
            15'd13913: data <= 8'h1F;
            15'd13914: data <= 8'h80;
            15'd13915: data <= 8'h00;
            15'd13916: data <= 8'h00;
            15'd13917: data <= 8'h00;
            15'd13918: data <= 8'h00;
            15'd13919: data <= 8'h00;
            15'd13920: data <= 8'h00;
            15'd13921: data <= 8'h00;
            15'd13922: data <= 8'h00;
            15'd13923: data <= 8'h00;
            15'd13924: data <= 8'h00;
            15'd13925: data <= 8'h03;
            15'd13926: data <= 8'hFF;
            15'd13927: data <= 8'hFF;
            15'd13928: data <= 8'hFF;
            15'd13929: data <= 8'hF8;
            15'd13930: data <= 8'h7E;
            15'd13931: data <= 8'h0F;
            15'd13932: data <= 8'hFF;
            15'd13933: data <= 8'hE0;
            15'd13934: data <= 8'h00;
            15'd13935: data <= 8'h00;
            15'd13936: data <= 8'h03;
            15'd13937: data <= 8'hFF;
            15'd13938: data <= 8'hFF;
            15'd13939: data <= 8'hFF;
            15'd13940: data <= 8'hFF;
            15'd13941: data <= 8'hFF;
            15'd13942: data <= 8'hE0;
            15'd13943: data <= 8'h1F;
            15'd13944: data <= 8'h80;
            15'd13945: data <= 8'h00;
            15'd13946: data <= 8'h00;
            15'd13947: data <= 8'h00;
            15'd13948: data <= 8'h00;
            15'd13949: data <= 8'h00;
            15'd13950: data <= 8'h00;
            15'd13951: data <= 8'h00;
            15'd13952: data <= 8'h00;
            15'd13953: data <= 8'h00;
            15'd13954: data <= 8'h00;
            15'd13955: data <= 8'h03;
            15'd13956: data <= 8'hFF;
            15'd13957: data <= 8'hFF;
            15'd13958: data <= 8'hFF;
            15'd13959: data <= 8'hF8;
            15'd13960: data <= 8'h7F;
            15'd13961: data <= 8'h0F;
            15'd13962: data <= 8'hFF;
            15'd13963: data <= 8'hF8;
            15'd13964: data <= 8'h00;
            15'd13965: data <= 8'h00;
            15'd13966: data <= 8'h07;
            15'd13967: data <= 8'hFF;
            15'd13968: data <= 8'hFF;
            15'd13969: data <= 8'hFF;
            15'd13970: data <= 8'hFF;
            15'd13971: data <= 8'hFF;
            15'd13972: data <= 8'hF0;
            15'd13973: data <= 8'h1F;
            15'd13974: data <= 8'h80;
            15'd13975: data <= 8'h00;
            15'd13976: data <= 8'h00;
            15'd13977: data <= 8'h00;
            15'd13978: data <= 8'h00;
            15'd13979: data <= 8'h00;
            15'd13980: data <= 8'h00;
            15'd13981: data <= 8'h00;
            15'd13982: data <= 8'h00;
            15'd13983: data <= 8'h00;
            15'd13984: data <= 8'h00;
            15'd13985: data <= 8'h03;
            15'd13986: data <= 8'hFF;
            15'd13987: data <= 8'hFF;
            15'd13988: data <= 8'hFF;
            15'd13989: data <= 8'hF8;
            15'd13990: data <= 8'h7F;
            15'd13991: data <= 8'h07;
            15'd13992: data <= 8'hFF;
            15'd13993: data <= 8'hFF;
            15'd13994: data <= 8'h00;
            15'd13995: data <= 8'h00;
            15'd13996: data <= 8'h1F;
            15'd13997: data <= 8'hFF;
            15'd13998: data <= 8'hFF;
            15'd13999: data <= 8'hFF;
            15'd14000: data <= 8'hFF;
            15'd14001: data <= 8'hFF;
            15'd14002: data <= 8'hF0;
            15'd14003: data <= 8'h1F;
            15'd14004: data <= 8'h80;
            15'd14005: data <= 8'h00;
            15'd14006: data <= 8'h00;
            15'd14007: data <= 8'h00;
            15'd14008: data <= 8'h00;
            15'd14009: data <= 8'h00;
            15'd14010: data <= 8'h00;
            15'd14011: data <= 8'h00;
            15'd14012: data <= 8'h00;
            15'd14013: data <= 8'h00;
            15'd14014: data <= 8'h00;
            15'd14015: data <= 8'h03;
            15'd14016: data <= 8'hFF;
            15'd14017: data <= 8'hFF;
            15'd14018: data <= 8'hFF;
            15'd14019: data <= 8'hF8;
            15'd14020: data <= 8'h7F;
            15'd14021: data <= 8'h87;
            15'd14022: data <= 8'hFF;
            15'd14023: data <= 8'hFF;
            15'd14024: data <= 8'hF0;
            15'd14025: data <= 8'h00;
            15'd14026: data <= 8'h7F;
            15'd14027: data <= 8'hFF;
            15'd14028: data <= 8'hFF;
            15'd14029: data <= 8'hFF;
            15'd14030: data <= 8'hFF;
            15'd14031: data <= 8'hFF;
            15'd14032: data <= 8'hF8;
            15'd14033: data <= 8'h0F;
            15'd14034: data <= 8'h80;
            15'd14035: data <= 8'h00;
            15'd14036: data <= 8'h00;
            15'd14037: data <= 8'h00;
            15'd14038: data <= 8'h00;
            15'd14039: data <= 8'h00;
            15'd14040: data <= 8'h00;
            15'd14041: data <= 8'h00;
            15'd14042: data <= 8'h00;
            15'd14043: data <= 8'h00;
            15'd14044: data <= 8'h00;
            15'd14045: data <= 8'h03;
            15'd14046: data <= 8'hFF;
            15'd14047: data <= 8'hFF;
            15'd14048: data <= 8'hFF;
            15'd14049: data <= 8'hF8;
            15'd14050: data <= 8'h7F;
            15'd14051: data <= 8'h83;
            15'd14052: data <= 8'hFF;
            15'd14053: data <= 8'hFF;
            15'd14054: data <= 8'hFE;
            15'd14055: data <= 8'h01;
            15'd14056: data <= 8'hFF;
            15'd14057: data <= 8'hFF;
            15'd14058: data <= 8'hFF;
            15'd14059: data <= 8'hFF;
            15'd14060: data <= 8'hFF;
            15'd14061: data <= 8'hFF;
            15'd14062: data <= 8'hF8;
            15'd14063: data <= 8'h0F;
            15'd14064: data <= 8'h80;
            15'd14065: data <= 8'h00;
            15'd14066: data <= 8'h00;
            15'd14067: data <= 8'h00;
            15'd14068: data <= 8'h00;
            15'd14069: data <= 8'h00;
            15'd14070: data <= 8'h00;
            15'd14071: data <= 8'h00;
            15'd14072: data <= 8'h00;
            15'd14073: data <= 8'h00;
            15'd14074: data <= 8'h00;
            15'd14075: data <= 8'h03;
            15'd14076: data <= 8'hFF;
            15'd14077: data <= 8'hFF;
            15'd14078: data <= 8'hFF;
            15'd14079: data <= 8'hF8;
            15'd14080: data <= 8'h7F;
            15'd14081: data <= 8'hC1;
            15'd14082: data <= 8'hFF;
            15'd14083: data <= 8'hFF;
            15'd14084: data <= 8'hFF;
            15'd14085: data <= 8'hFF;
            15'd14086: data <= 8'hFF;
            15'd14087: data <= 8'hFF;
            15'd14088: data <= 8'hFF;
            15'd14089: data <= 8'hFF;
            15'd14090: data <= 8'hFF;
            15'd14091: data <= 8'hFF;
            15'd14092: data <= 8'hF8;
            15'd14093: data <= 8'h0F;
            15'd14094: data <= 8'h80;
            15'd14095: data <= 8'h00;
            15'd14096: data <= 8'h00;
            15'd14097: data <= 8'h00;
            15'd14098: data <= 8'h00;
            15'd14099: data <= 8'h00;
            15'd14100: data <= 8'h00;
            15'd14101: data <= 8'h00;
            15'd14102: data <= 8'h00;
            15'd14103: data <= 8'h00;
            15'd14104: data <= 8'h00;
            15'd14105: data <= 8'h03;
            15'd14106: data <= 8'hFF;
            15'd14107: data <= 8'hFF;
            15'd14108: data <= 8'hFF;
            15'd14109: data <= 8'hF8;
            15'd14110: data <= 8'h7F;
            15'd14111: data <= 8'hC1;
            15'd14112: data <= 8'hFF;
            15'd14113: data <= 8'hFF;
            15'd14114: data <= 8'hFF;
            15'd14115: data <= 8'hFF;
            15'd14116: data <= 8'hFF;
            15'd14117: data <= 8'hFF;
            15'd14118: data <= 8'hFF;
            15'd14119: data <= 8'hFF;
            15'd14120: data <= 8'hFF;
            15'd14121: data <= 8'hFF;
            15'd14122: data <= 8'hF8;
            15'd14123: data <= 8'h07;
            15'd14124: data <= 8'h80;
            15'd14125: data <= 8'h00;
            15'd14126: data <= 8'h00;
            15'd14127: data <= 8'h00;
            15'd14128: data <= 8'h00;
            15'd14129: data <= 8'h00;
            15'd14130: data <= 8'h00;
            15'd14131: data <= 8'h00;
            15'd14132: data <= 8'h00;
            15'd14133: data <= 8'h00;
            15'd14134: data <= 8'h00;
            15'd14135: data <= 8'h03;
            15'd14136: data <= 8'hFF;
            15'd14137: data <= 8'hFF;
            15'd14138: data <= 8'hFF;
            15'd14139: data <= 8'hF8;
            15'd14140: data <= 8'h7F;
            15'd14141: data <= 8'hE0;
            15'd14142: data <= 8'hFF;
            15'd14143: data <= 8'hFF;
            15'd14144: data <= 8'hFF;
            15'd14145: data <= 8'hFF;
            15'd14146: data <= 8'hFF;
            15'd14147: data <= 8'hFF;
            15'd14148: data <= 8'hFF;
            15'd14149: data <= 8'hFF;
            15'd14150: data <= 8'hFF;
            15'd14151: data <= 8'hFF;
            15'd14152: data <= 8'hFC;
            15'd14153: data <= 8'h07;
            15'd14154: data <= 8'h80;
            15'd14155: data <= 8'h00;
            15'd14156: data <= 8'h00;
            15'd14157: data <= 8'h00;
            15'd14158: data <= 8'h00;
            15'd14159: data <= 8'h00;
            15'd14160: data <= 8'h00;
            15'd14161: data <= 8'h00;
            15'd14162: data <= 8'h00;
            15'd14163: data <= 8'h00;
            15'd14164: data <= 8'h00;
            15'd14165: data <= 8'h03;
            15'd14166: data <= 8'hFF;
            15'd14167: data <= 8'hFF;
            15'd14168: data <= 8'hFF;
            15'd14169: data <= 8'hFC;
            15'd14170: data <= 8'h7F;
            15'd14171: data <= 8'hE0;
            15'd14172: data <= 8'h7F;
            15'd14173: data <= 8'hFF;
            15'd14174: data <= 8'hFF;
            15'd14175: data <= 8'hFF;
            15'd14176: data <= 8'hFF;
            15'd14177: data <= 8'hFF;
            15'd14178: data <= 8'hFF;
            15'd14179: data <= 8'hFF;
            15'd14180: data <= 8'hFF;
            15'd14181: data <= 8'hFF;
            15'd14182: data <= 8'hFC;
            15'd14183: data <= 8'h07;
            15'd14184: data <= 8'h80;
            15'd14185: data <= 8'h00;
            15'd14186: data <= 8'h00;
            15'd14187: data <= 8'h00;
            15'd14188: data <= 8'h00;
            15'd14189: data <= 8'h00;
            15'd14190: data <= 8'h00;
            15'd14191: data <= 8'h00;
            15'd14192: data <= 8'h00;
            15'd14193: data <= 8'h00;
            15'd14194: data <= 8'h00;
            15'd14195: data <= 8'h03;
            15'd14196: data <= 8'hFF;
            15'd14197: data <= 8'hFF;
            15'd14198: data <= 8'hFF;
            15'd14199: data <= 8'hFC;
            15'd14200: data <= 8'h7F;
            15'd14201: data <= 8'hF0;
            15'd14202: data <= 8'h7F;
            15'd14203: data <= 8'hFF;
            15'd14204: data <= 8'hFF;
            15'd14205: data <= 8'hFF;
            15'd14206: data <= 8'hFF;
            15'd14207: data <= 8'hFF;
            15'd14208: data <= 8'hFF;
            15'd14209: data <= 8'hFF;
            15'd14210: data <= 8'hFF;
            15'd14211: data <= 8'hFF;
            15'd14212: data <= 8'hFC;
            15'd14213: data <= 8'h03;
            15'd14214: data <= 8'h80;
            15'd14215: data <= 8'h00;
            15'd14216: data <= 8'h00;
            15'd14217: data <= 8'h00;
            15'd14218: data <= 8'h00;
            15'd14219: data <= 8'h00;
            15'd14220: data <= 8'h00;
            15'd14221: data <= 8'h00;
            15'd14222: data <= 8'h00;
            15'd14223: data <= 8'h00;
            15'd14224: data <= 8'h00;
            15'd14225: data <= 8'h03;
            15'd14226: data <= 8'hFF;
            15'd14227: data <= 8'hFF;
            15'd14228: data <= 8'hFF;
            15'd14229: data <= 8'hFC;
            15'd14230: data <= 8'h7F;
            15'd14231: data <= 8'hF8;
            15'd14232: data <= 8'h3F;
            15'd14233: data <= 8'hFF;
            15'd14234: data <= 8'hFF;
            15'd14235: data <= 8'hFF;
            15'd14236: data <= 8'hFF;
            15'd14237: data <= 8'hFF;
            15'd14238: data <= 8'hFF;
            15'd14239: data <= 8'hFF;
            15'd14240: data <= 8'hFF;
            15'd14241: data <= 8'hFF;
            15'd14242: data <= 8'hFE;
            15'd14243: data <= 8'h03;
            15'd14244: data <= 8'h80;
            15'd14245: data <= 8'h00;
            15'd14246: data <= 8'h00;
            15'd14247: data <= 8'h00;
            15'd14248: data <= 8'h00;
            15'd14249: data <= 8'h00;
            15'd14250: data <= 8'h00;
            15'd14251: data <= 8'h00;
            15'd14252: data <= 8'h00;
            15'd14253: data <= 8'h00;
            15'd14254: data <= 8'h00;
            15'd14255: data <= 8'h03;
            15'd14256: data <= 8'hFF;
            15'd14257: data <= 8'hFF;
            15'd14258: data <= 8'hFF;
            15'd14259: data <= 8'hFC;
            15'd14260: data <= 8'h7F;
            15'd14261: data <= 8'hFC;
            15'd14262: data <= 8'h1F;
            15'd14263: data <= 8'hFF;
            15'd14264: data <= 8'hFF;
            15'd14265: data <= 8'hFF;
            15'd14266: data <= 8'hFF;
            15'd14267: data <= 8'hFF;
            15'd14268: data <= 8'hFF;
            15'd14269: data <= 8'hFF;
            15'd14270: data <= 8'hFF;
            15'd14271: data <= 8'hFF;
            15'd14272: data <= 8'hFE;
            15'd14273: data <= 8'h03;
            15'd14274: data <= 8'h80;
            15'd14275: data <= 8'h00;
            15'd14276: data <= 8'h00;
            15'd14277: data <= 8'h00;
            15'd14278: data <= 8'h00;
            15'd14279: data <= 8'h00;
            15'd14280: data <= 8'h00;
            15'd14281: data <= 8'h00;
            15'd14282: data <= 8'h00;
            15'd14283: data <= 8'h00;
            15'd14284: data <= 8'h00;
            15'd14285: data <= 8'h03;
            15'd14286: data <= 8'hFF;
            15'd14287: data <= 8'hFF;
            15'd14288: data <= 8'hFF;
            15'd14289: data <= 8'hFC;
            15'd14290: data <= 8'h7F;
            15'd14291: data <= 8'hFC;
            15'd14292: data <= 8'h0F;
            15'd14293: data <= 8'hFF;
            15'd14294: data <= 8'hFF;
            15'd14295: data <= 8'hFF;
            15'd14296: data <= 8'hFF;
            15'd14297: data <= 8'hFF;
            15'd14298: data <= 8'hFF;
            15'd14299: data <= 8'hFF;
            15'd14300: data <= 8'hFF;
            15'd14301: data <= 8'hFF;
            15'd14302: data <= 8'hFE;
            15'd14303: data <= 8'h03;
            15'd14304: data <= 8'h80;
            15'd14305: data <= 8'h00;
            15'd14306: data <= 8'h00;
            15'd14307: data <= 8'h00;
            15'd14308: data <= 8'h00;
            15'd14309: data <= 8'h00;
            15'd14310: data <= 8'h00;
            15'd14311: data <= 8'h00;
            15'd14312: data <= 8'h00;
            15'd14313: data <= 8'h00;
            15'd14314: data <= 8'h00;
            15'd14315: data <= 8'h03;
            15'd14316: data <= 8'hFF;
            15'd14317: data <= 8'hFF;
            15'd14318: data <= 8'hFF;
            15'd14319: data <= 8'hFC;
            15'd14320: data <= 8'h7F;
            15'd14321: data <= 8'hFE;
            15'd14322: data <= 8'h07;
            15'd14323: data <= 8'hFF;
            15'd14324: data <= 8'hFF;
            15'd14325: data <= 8'hFF;
            15'd14326: data <= 8'hFF;
            15'd14327: data <= 8'hFF;
            15'd14328: data <= 8'hFF;
            15'd14329: data <= 8'hFF;
            15'd14330: data <= 8'hFF;
            15'd14331: data <= 8'hFF;
            15'd14332: data <= 8'hFF;
            15'd14333: data <= 8'h03;
            15'd14334: data <= 8'h80;
            15'd14335: data <= 8'h00;
            15'd14336: data <= 8'h00;
            15'd14337: data <= 8'h00;
            15'd14338: data <= 8'h00;
            15'd14339: data <= 8'h00;
            15'd14340: data <= 8'h00;
            15'd14341: data <= 8'h00;
            15'd14342: data <= 8'h00;
            15'd14343: data <= 8'h00;
            15'd14344: data <= 8'h00;
            15'd14345: data <= 8'h03;
            15'd14346: data <= 8'hFF;
            15'd14347: data <= 8'hFF;
            15'd14348: data <= 8'hFF;
            15'd14349: data <= 8'hFC;
            15'd14350: data <= 8'h7F;
            15'd14351: data <= 8'hFF;
            15'd14352: data <= 8'h03;
            15'd14353: data <= 8'hFF;
            15'd14354: data <= 8'hFF;
            15'd14355: data <= 8'hFF;
            15'd14356: data <= 8'hFF;
            15'd14357: data <= 8'hFF;
            15'd14358: data <= 8'hFF;
            15'd14359: data <= 8'hFF;
            15'd14360: data <= 8'hFF;
            15'd14361: data <= 8'hFF;
            15'd14362: data <= 8'hFF;
            15'd14363: data <= 8'h01;
            15'd14364: data <= 8'h80;
            15'd14365: data <= 8'h00;
            15'd14366: data <= 8'h00;
            15'd14367: data <= 8'h00;
            15'd14368: data <= 8'h00;
            15'd14369: data <= 8'h00;
            15'd14370: data <= 8'h00;
            15'd14371: data <= 8'h00;
            15'd14372: data <= 8'h00;
            15'd14373: data <= 8'h00;
            15'd14374: data <= 8'h00;
            15'd14375: data <= 8'h03;
            15'd14376: data <= 8'hFF;
            15'd14377: data <= 8'hFF;
            15'd14378: data <= 8'hFF;
            15'd14379: data <= 8'hFC;
            15'd14380: data <= 8'h7F;
            15'd14381: data <= 8'hFF;
            15'd14382: data <= 8'h81;
            15'd14383: data <= 8'hFF;
            15'd14384: data <= 8'hFF;
            15'd14385: data <= 8'hFF;
            15'd14386: data <= 8'hFF;
            15'd14387: data <= 8'hFF;
            15'd14388: data <= 8'hFF;
            15'd14389: data <= 8'hFF;
            15'd14390: data <= 8'hFF;
            15'd14391: data <= 8'hFF;
            15'd14392: data <= 8'hFF;
            15'd14393: data <= 8'h81;
            15'd14394: data <= 8'h80;
            15'd14395: data <= 8'h00;
            15'd14396: data <= 8'h00;
            15'd14397: data <= 8'h00;
            15'd14398: data <= 8'h00;
            15'd14399: data <= 8'h00;
            15'd14400: data <= 8'h00;
            15'd14401: data <= 8'h00;
            15'd14402: data <= 8'h00;
            15'd14403: data <= 8'h00;
            15'd14404: data <= 8'h00;
            15'd14405: data <= 8'h03;
            15'd14406: data <= 8'hFF;
            15'd14407: data <= 8'hFF;
            15'd14408: data <= 8'hFF;
            15'd14409: data <= 8'hFC;
            15'd14410: data <= 8'h7F;
            15'd14411: data <= 8'hFF;
            15'd14412: data <= 8'hC1;
            15'd14413: data <= 8'hFF;
            15'd14414: data <= 8'hFF;
            15'd14415: data <= 8'hFF;
            15'd14416: data <= 8'hFF;
            15'd14417: data <= 8'hFF;
            15'd14418: data <= 8'hFF;
            15'd14419: data <= 8'hFF;
            15'd14420: data <= 8'hFF;
            15'd14421: data <= 8'hFF;
            15'd14422: data <= 8'hFF;
            15'd14423: data <= 8'h81;
            15'd14424: data <= 8'h80;
            15'd14425: data <= 8'h00;
            15'd14426: data <= 8'h00;
            15'd14427: data <= 8'h00;
            15'd14428: data <= 8'h00;
            15'd14429: data <= 8'h00;
            15'd14430: data <= 8'h00;
            15'd14431: data <= 8'h00;
            15'd14432: data <= 8'h00;
            15'd14433: data <= 8'h00;
            15'd14434: data <= 8'h00;
            15'd14435: data <= 8'h03;
            15'd14436: data <= 8'hFF;
            15'd14437: data <= 8'hFF;
            15'd14438: data <= 8'hFF;
            15'd14439: data <= 8'hF8;
            15'd14440: data <= 8'h7F;
            15'd14441: data <= 8'hFF;
            15'd14442: data <= 8'hE0;
            15'd14443: data <= 8'h7F;
            15'd14444: data <= 8'hFF;
            15'd14445: data <= 8'hFF;
            15'd14446: data <= 8'hFF;
            15'd14447: data <= 8'hFF;
            15'd14448: data <= 8'hFF;
            15'd14449: data <= 8'hFF;
            15'd14450: data <= 8'hFF;
            15'd14451: data <= 8'hFF;
            15'd14452: data <= 8'hFF;
            15'd14453: data <= 8'h81;
            15'd14454: data <= 8'h80;
            15'd14455: data <= 8'h00;
            15'd14456: data <= 8'h00;
            15'd14457: data <= 8'h00;
            15'd14458: data <= 8'h00;
            15'd14459: data <= 8'h00;
            15'd14460: data <= 8'h00;
            15'd14461: data <= 8'h00;
            15'd14462: data <= 8'h00;
            15'd14463: data <= 8'h00;
            15'd14464: data <= 8'h00;
            15'd14465: data <= 8'h03;
            15'd14466: data <= 8'hFF;
            15'd14467: data <= 8'hFF;
            15'd14468: data <= 8'hFF;
            15'd14469: data <= 8'hF0;
            15'd14470: data <= 8'h7F;
            15'd14471: data <= 8'hFF;
            15'd14472: data <= 8'hF0;
            15'd14473: data <= 8'h3F;
            15'd14474: data <= 8'hFF;
            15'd14475: data <= 8'hFF;
            15'd14476: data <= 8'hFF;
            15'd14477: data <= 8'hFF;
            15'd14478: data <= 8'hFF;
            15'd14479: data <= 8'hFF;
            15'd14480: data <= 8'hFF;
            15'd14481: data <= 8'hFF;
            15'd14482: data <= 8'hFF;
            15'd14483: data <= 8'h80;
            15'd14484: data <= 8'h80;
            15'd14485: data <= 8'h00;
            15'd14486: data <= 8'h00;
            15'd14487: data <= 8'h00;
            15'd14488: data <= 8'h00;
            15'd14489: data <= 8'h00;
            15'd14490: data <= 8'h00;
            15'd14491: data <= 8'h00;
            15'd14492: data <= 8'h00;
            15'd14493: data <= 8'h00;
            15'd14494: data <= 8'h00;
            15'd14495: data <= 8'h03;
            15'd14496: data <= 8'hFF;
            15'd14497: data <= 8'hFF;
            15'd14498: data <= 8'hFF;
            15'd14499: data <= 8'hF0;
            15'd14500: data <= 8'h7F;
            15'd14501: data <= 8'hFF;
            15'd14502: data <= 8'hF0;
            15'd14503: data <= 8'h1F;
            15'd14504: data <= 8'hFF;
            15'd14505: data <= 8'hFF;
            15'd14506: data <= 8'hFF;
            15'd14507: data <= 8'hFF;
            15'd14508: data <= 8'hFF;
            15'd14509: data <= 8'hFF;
            15'd14510: data <= 8'hFF;
            15'd14511: data <= 8'hFF;
            15'd14512: data <= 8'hFF;
            15'd14513: data <= 8'h80;
            15'd14514: data <= 8'h80;
            15'd14515: data <= 8'h00;
            15'd14516: data <= 8'h00;
            15'd14517: data <= 8'h00;
            15'd14518: data <= 8'h00;
            15'd14519: data <= 8'h00;
            15'd14520: data <= 8'h00;
            15'd14521: data <= 8'h00;
            15'd14522: data <= 8'h00;
            15'd14523: data <= 8'h00;
            15'd14524: data <= 8'h00;
            15'd14525: data <= 8'h03;
            15'd14526: data <= 8'hFF;
            15'd14527: data <= 8'hFF;
            15'd14528: data <= 8'hFF;
            15'd14529: data <= 8'hF0;
            15'd14530: data <= 8'h3F;
            15'd14531: data <= 8'hFF;
            15'd14532: data <= 8'hF8;
            15'd14533: data <= 8'h07;
            15'd14534: data <= 8'hFF;
            15'd14535: data <= 8'hFF;
            15'd14536: data <= 8'hFF;
            15'd14537: data <= 8'hFF;
            15'd14538: data <= 8'hFF;
            15'd14539: data <= 8'hFF;
            15'd14540: data <= 8'hFF;
            15'd14541: data <= 8'hFF;
            15'd14542: data <= 8'hFF;
            15'd14543: data <= 8'h80;
            15'd14544: data <= 8'h80;
            15'd14545: data <= 8'h00;
            15'd14546: data <= 8'h00;
            15'd14547: data <= 8'h00;
            15'd14548: data <= 8'h00;
            15'd14549: data <= 8'h00;
            15'd14550: data <= 8'h00;
            15'd14551: data <= 8'h00;
            15'd14552: data <= 8'h00;
            15'd14553: data <= 8'h00;
            15'd14554: data <= 8'h00;
            15'd14555: data <= 8'h03;
            15'd14556: data <= 8'hFF;
            15'd14557: data <= 8'hFF;
            15'd14558: data <= 8'hFF;
            15'd14559: data <= 8'hF8;
            15'd14560: data <= 8'h3F;
            15'd14561: data <= 8'hFF;
            15'd14562: data <= 8'hFE;
            15'd14563: data <= 8'h01;
            15'd14564: data <= 8'hFF;
            15'd14565: data <= 8'hFF;
            15'd14566: data <= 8'hFF;
            15'd14567: data <= 8'hFF;
            15'd14568: data <= 8'hFF;
            15'd14569: data <= 8'hFF;
            15'd14570: data <= 8'hFF;
            15'd14571: data <= 8'hFF;
            15'd14572: data <= 8'hFF;
            15'd14573: data <= 8'hC0;
            15'd14574: data <= 8'h00;
            15'd14575: data <= 8'h00;
            15'd14576: data <= 8'h00;
            15'd14577: data <= 8'h00;
            15'd14578: data <= 8'h00;
            15'd14579: data <= 8'h00;
            15'd14580: data <= 8'h00;
            15'd14581: data <= 8'h00;
            15'd14582: data <= 8'h00;
            15'd14583: data <= 8'h00;
            15'd14584: data <= 8'h00;
            15'd14585: data <= 8'h03;
            15'd14586: data <= 8'hFF;
            15'd14587: data <= 8'hFF;
            15'd14588: data <= 8'hFF;
            15'd14589: data <= 8'hF8;
            15'd14590: data <= 8'h3F;
            15'd14591: data <= 8'hFF;
            15'd14592: data <= 8'hFF;
            15'd14593: data <= 8'h00;
            15'd14594: data <= 8'hFF;
            15'd14595: data <= 8'hFF;
            15'd14596: data <= 8'hFF;
            15'd14597: data <= 8'hFF;
            15'd14598: data <= 8'hFF;
            15'd14599: data <= 8'hFF;
            15'd14600: data <= 8'hFF;
            15'd14601: data <= 8'hFF;
            15'd14602: data <= 8'hFF;
            15'd14603: data <= 8'hC0;
            15'd14604: data <= 8'h00;
            15'd14605: data <= 8'h00;
            15'd14606: data <= 8'h00;
            15'd14607: data <= 8'h00;
            15'd14608: data <= 8'h00;
            15'd14609: data <= 8'h00;
            15'd14610: data <= 8'h00;
            15'd14611: data <= 8'h00;
            15'd14612: data <= 8'h00;
            15'd14613: data <= 8'h00;
            15'd14614: data <= 8'h00;
            15'd14615: data <= 8'h03;
            15'd14616: data <= 8'hFF;
            15'd14617: data <= 8'hFF;
            15'd14618: data <= 8'hFF;
            15'd14619: data <= 8'hF8;
            15'd14620: data <= 8'h7F;
            15'd14621: data <= 8'hFF;
            15'd14622: data <= 8'hFF;
            15'd14623: data <= 8'h80;
            15'd14624: data <= 8'h1F;
            15'd14625: data <= 8'hFF;
            15'd14626: data <= 8'hFF;
            15'd14627: data <= 8'hFF;
            15'd14628: data <= 8'hFF;
            15'd14629: data <= 8'hFF;
            15'd14630: data <= 8'hFF;
            15'd14631: data <= 8'hFF;
            15'd14632: data <= 8'hFF;
            15'd14633: data <= 8'hC0;
            15'd14634: data <= 8'h00;
            15'd14635: data <= 8'h00;
            15'd14636: data <= 8'h00;
            15'd14637: data <= 8'h00;
            15'd14638: data <= 8'h00;
            15'd14639: data <= 8'h00;
            15'd14640: data <= 8'h00;
            15'd14641: data <= 8'h00;
            15'd14642: data <= 8'h00;
            15'd14643: data <= 8'h00;
            15'd14644: data <= 8'h00;
            15'd14645: data <= 8'h03;
            15'd14646: data <= 8'hFF;
            15'd14647: data <= 8'hFF;
            15'd14648: data <= 8'hFF;
            15'd14649: data <= 8'hF8;
            15'd14650: data <= 8'h7F;
            15'd14651: data <= 8'hFF;
            15'd14652: data <= 8'hFF;
            15'd14653: data <= 8'hC0;
            15'd14654: data <= 8'h07;
            15'd14655: data <= 8'hFF;
            15'd14656: data <= 8'hFF;
            15'd14657: data <= 8'hFF;
            15'd14658: data <= 8'hFF;
            15'd14659: data <= 8'hFF;
            15'd14660: data <= 8'hFF;
            15'd14661: data <= 8'hFF;
            15'd14662: data <= 8'hFF;
            15'd14663: data <= 8'hC0;
            15'd14664: data <= 8'h00;
            15'd14665: data <= 8'h00;
            15'd14666: data <= 8'h00;
            15'd14667: data <= 8'h00;
            15'd14668: data <= 8'h00;
            15'd14669: data <= 8'h00;
            15'd14670: data <= 8'h00;
            15'd14671: data <= 8'h00;
            15'd14672: data <= 8'h00;
            15'd14673: data <= 8'h00;
            15'd14674: data <= 8'h00;
            15'd14675: data <= 8'h03;
            15'd14676: data <= 8'hFF;
            15'd14677: data <= 8'hFF;
            15'd14678: data <= 8'hFF;
            15'd14679: data <= 8'hF8;
            15'd14680: data <= 8'h7F;
            15'd14681: data <= 8'hFF;
            15'd14682: data <= 8'hFF;
            15'd14683: data <= 8'hE0;
            15'd14684: data <= 8'h01;
            15'd14685: data <= 8'hFF;
            15'd14686: data <= 8'hFF;
            15'd14687: data <= 8'hFF;
            15'd14688: data <= 8'hFF;
            15'd14689: data <= 8'hFF;
            15'd14690: data <= 8'hFF;
            15'd14691: data <= 8'hFF;
            15'd14692: data <= 8'hFF;
            15'd14693: data <= 8'hC0;
            15'd14694: data <= 8'h00;
            15'd14695: data <= 8'h00;
            15'd14696: data <= 8'h00;
            15'd14697: data <= 8'h00;
            15'd14698: data <= 8'h00;
            15'd14699: data <= 8'h00;
            15'd14700: data <= 8'h00;
            15'd14701: data <= 8'h00;
            15'd14702: data <= 8'h00;
            15'd14703: data <= 8'h00;
            15'd14704: data <= 8'h00;
            15'd14705: data <= 8'h03;
            15'd14706: data <= 8'hFF;
            15'd14707: data <= 8'hFF;
            15'd14708: data <= 8'hFF;
            15'd14709: data <= 8'hF8;
            15'd14710: data <= 8'h7F;
            15'd14711: data <= 8'hFF;
            15'd14712: data <= 8'hFF;
            15'd14713: data <= 8'hF8;
            15'd14714: data <= 8'h00;
            15'd14715: data <= 8'h7F;
            15'd14716: data <= 8'hFC;
            15'd14717: data <= 8'h7F;
            15'd14718: data <= 8'hFF;
            15'd14719: data <= 8'hFF;
            15'd14720: data <= 8'hFF;
            15'd14721: data <= 8'hFF;
            15'd14722: data <= 8'hFF;
            15'd14723: data <= 8'hE0;
            15'd14724: data <= 8'h00;
            15'd14725: data <= 8'h00;
            15'd14726: data <= 8'h00;
            15'd14727: data <= 8'h00;
            15'd14728: data <= 8'h00;
            15'd14729: data <= 8'h00;
            15'd14730: data <= 8'h00;
            15'd14731: data <= 8'h00;
            15'd14732: data <= 8'h00;
            15'd14733: data <= 8'h00;
            15'd14734: data <= 8'h00;
            15'd14735: data <= 8'h03;
            15'd14736: data <= 8'hFF;
            15'd14737: data <= 8'hFF;
            15'd14738: data <= 8'hFF;
            15'd14739: data <= 8'hF8;
            15'd14740: data <= 8'h7F;
            15'd14741: data <= 8'hFF;
            15'd14742: data <= 8'hFF;
            15'd14743: data <= 8'hFC;
            15'd14744: data <= 8'h00;
            15'd14745: data <= 8'h00;
            15'd14746: data <= 8'hC0;
            15'd14747: data <= 8'h3F;
            15'd14748: data <= 8'hFF;
            15'd14749: data <= 8'hFF;
            15'd14750: data <= 8'hFF;
            15'd14751: data <= 8'hFF;
            15'd14752: data <= 8'hFF;
            15'd14753: data <= 8'hE0;
            15'd14754: data <= 8'h00;
            15'd14755: data <= 8'h00;
            15'd14756: data <= 8'h00;
            15'd14757: data <= 8'h00;
            15'd14758: data <= 8'h00;
            15'd14759: data <= 8'h00;
            15'd14760: data <= 8'h00;
            15'd14761: data <= 8'h00;
            15'd14762: data <= 8'h00;
            15'd14763: data <= 8'h00;
            15'd14764: data <= 8'h00;
            15'd14765: data <= 8'h03;
            15'd14766: data <= 8'hFF;
            15'd14767: data <= 8'hFF;
            15'd14768: data <= 8'hFF;
            15'd14769: data <= 8'hF0;
            15'd14770: data <= 8'h7F;
            15'd14771: data <= 8'hFF;
            15'd14772: data <= 8'hFF;
            15'd14773: data <= 8'hFF;
            15'd14774: data <= 8'h00;
            15'd14775: data <= 8'h00;
            15'd14776: data <= 8'h00;
            15'd14777: data <= 8'h1F;
            15'd14778: data <= 8'hFF;
            15'd14779: data <= 8'hFF;
            15'd14780: data <= 8'hFF;
            15'd14781: data <= 8'hFF;
            15'd14782: data <= 8'hFF;
            15'd14783: data <= 8'hE0;
            15'd14784: data <= 8'h00;
            15'd14785: data <= 8'h00;
            15'd14786: data <= 8'h00;
            15'd14787: data <= 8'h00;
            15'd14788: data <= 8'h00;
            15'd14789: data <= 8'h00;
            15'd14790: data <= 8'h00;
            15'd14791: data <= 8'h00;
            15'd14792: data <= 8'h00;
            15'd14793: data <= 8'h00;
            15'd14794: data <= 8'h00;
            15'd14795: data <= 8'h03;
            15'd14796: data <= 8'hFF;
            15'd14797: data <= 8'hFF;
            15'd14798: data <= 8'hFF;
            15'd14799: data <= 8'hF0;
            15'd14800: data <= 8'h7F;
            15'd14801: data <= 8'hFF;
            15'd14802: data <= 8'hFF;
            15'd14803: data <= 8'hFF;
            15'd14804: data <= 8'hC0;
            15'd14805: data <= 8'h00;
            15'd14806: data <= 8'h00;
            15'd14807: data <= 8'h3F;
            15'd14808: data <= 8'hFF;
            15'd14809: data <= 8'hFF;
            15'd14810: data <= 8'hFF;
            15'd14811: data <= 8'hFF;
            15'd14812: data <= 8'hFF;
            15'd14813: data <= 8'hE0;
            15'd14814: data <= 8'h00;
            15'd14815: data <= 8'h00;
            15'd14816: data <= 8'h00;
            15'd14817: data <= 8'h00;
            15'd14818: data <= 8'h00;
            15'd14819: data <= 8'h00;
            15'd14820: data <= 8'h00;
            15'd14821: data <= 8'h00;
            15'd14822: data <= 8'h00;
            15'd14823: data <= 8'h00;
            15'd14824: data <= 8'h00;
            15'd14825: data <= 8'h03;
            15'd14826: data <= 8'hFF;
            15'd14827: data <= 8'hFF;
            15'd14828: data <= 8'hFF;
            15'd14829: data <= 8'hF0;
            15'd14830: data <= 8'h7F;
            15'd14831: data <= 8'hFF;
            15'd14832: data <= 8'hFF;
            15'd14833: data <= 8'hFF;
            15'd14834: data <= 8'hF0;
            15'd14835: data <= 8'h00;
            15'd14836: data <= 8'h00;
            15'd14837: data <= 8'h3F;
            15'd14838: data <= 8'hFF;
            15'd14839: data <= 8'hFF;
            15'd14840: data <= 8'hFF;
            15'd14841: data <= 8'hFF;
            15'd14842: data <= 8'hFF;
            15'd14843: data <= 8'hE0;
            15'd14844: data <= 8'h00;
            15'd14845: data <= 8'h00;
            15'd14846: data <= 8'h00;
            15'd14847: data <= 8'h00;
            15'd14848: data <= 8'h00;
            15'd14849: data <= 8'h00;
            15'd14850: data <= 8'h00;
            15'd14851: data <= 8'h00;
            15'd14852: data <= 8'h00;
            15'd14853: data <= 8'h00;
            15'd14854: data <= 8'h00;
            15'd14855: data <= 8'h03;
            15'd14856: data <= 8'hFF;
            15'd14857: data <= 8'hFF;
            15'd14858: data <= 8'hFF;
            15'd14859: data <= 8'hF0;
            15'd14860: data <= 8'h7F;
            15'd14861: data <= 8'hFF;
            15'd14862: data <= 8'hFF;
            15'd14863: data <= 8'hFF;
            15'd14864: data <= 8'hF8;
            15'd14865: data <= 8'h00;
            15'd14866: data <= 8'h00;
            15'd14867: data <= 8'h7F;
            15'd14868: data <= 8'hFF;
            15'd14869: data <= 8'hFF;
            15'd14870: data <= 8'hFF;
            15'd14871: data <= 8'hFF;
            15'd14872: data <= 8'hFF;
            15'd14873: data <= 8'hE0;
            15'd14874: data <= 8'h00;
            15'd14875: data <= 8'h00;
            15'd14876: data <= 8'h00;
            15'd14877: data <= 8'h00;
            15'd14878: data <= 8'h00;
            15'd14879: data <= 8'h00;
            15'd14880: data <= 8'h00;
            15'd14881: data <= 8'h00;
            15'd14882: data <= 8'h00;
            15'd14883: data <= 8'h00;
            15'd14884: data <= 8'h00;
            15'd14885: data <= 8'h03;
            15'd14886: data <= 8'hFF;
            15'd14887: data <= 8'hFF;
            15'd14888: data <= 8'hFF;
            15'd14889: data <= 8'hF0;
            15'd14890: data <= 8'h7F;
            15'd14891: data <= 8'hFF;
            15'd14892: data <= 8'hFF;
            15'd14893: data <= 8'hFF;
            15'd14894: data <= 8'hFF;
            15'd14895: data <= 8'hC0;
            15'd14896: data <= 8'h03;
            15'd14897: data <= 8'hFF;
            15'd14898: data <= 8'hFF;
            15'd14899: data <= 8'hFF;
            15'd14900: data <= 8'hFF;
            15'd14901: data <= 8'hFF;
            15'd14902: data <= 8'hFF;
            15'd14903: data <= 8'hF0;
            15'd14904: data <= 8'h00;
            15'd14905: data <= 8'h00;
            15'd14906: data <= 8'h00;
            15'd14907: data <= 8'h00;
            15'd14908: data <= 8'h00;
            15'd14909: data <= 8'h00;
            15'd14910: data <= 8'h00;
            15'd14911: data <= 8'h00;
            15'd14912: data <= 8'h00;
            15'd14913: data <= 8'h00;
            15'd14914: data <= 8'h00;
            15'd14915: data <= 8'h03;
            15'd14916: data <= 8'hFF;
            15'd14917: data <= 8'hFF;
            15'd14918: data <= 8'hFF;
            15'd14919: data <= 8'hF0;
            15'd14920: data <= 8'h7F;
            15'd14921: data <= 8'hFF;
            15'd14922: data <= 8'hFF;
            15'd14923: data <= 8'hFF;
            15'd14924: data <= 8'hFF;
            15'd14925: data <= 8'hFF;
            15'd14926: data <= 8'hFF;
            15'd14927: data <= 8'hFF;
            15'd14928: data <= 8'hFF;
            15'd14929: data <= 8'hFF;
            15'd14930: data <= 8'hFF;
            15'd14931: data <= 8'hFF;
            15'd14932: data <= 8'hFF;
            15'd14933: data <= 8'hF0;
            15'd14934: data <= 8'h00;
            15'd14935: data <= 8'h00;
            15'd14936: data <= 8'h00;
            15'd14937: data <= 8'h00;
            15'd14938: data <= 8'h00;
            15'd14939: data <= 8'h00;
            15'd14940: data <= 8'h00;
            15'd14941: data <= 8'h00;
            15'd14942: data <= 8'h00;
            15'd14943: data <= 8'h00;
            15'd14944: data <= 8'h00;
            15'd14945: data <= 8'h03;
            15'd14946: data <= 8'hFF;
            15'd14947: data <= 8'hFF;
            15'd14948: data <= 8'hFF;
            15'd14949: data <= 8'hF0;
            15'd14950: data <= 8'h7F;
            15'd14951: data <= 8'hFF;
            15'd14952: data <= 8'hFF;
            15'd14953: data <= 8'hFF;
            15'd14954: data <= 8'hFF;
            15'd14955: data <= 8'hFF;
            15'd14956: data <= 8'hFF;
            15'd14957: data <= 8'hFF;
            15'd14958: data <= 8'hFF;
            15'd14959: data <= 8'hFF;
            15'd14960: data <= 8'hFF;
            15'd14961: data <= 8'hFF;
            15'd14962: data <= 8'hFF;
            15'd14963: data <= 8'hF0;
            15'd14964: data <= 8'h00;
            15'd14965: data <= 8'h00;
            15'd14966: data <= 8'h00;
            15'd14967: data <= 8'h00;
            15'd14968: data <= 8'h00;
            15'd14969: data <= 8'h00;
            15'd14970: data <= 8'h00;
            15'd14971: data <= 8'h00;
            15'd14972: data <= 8'h00;
            15'd14973: data <= 8'h00;
            15'd14974: data <= 8'h00;
            15'd14975: data <= 8'h03;
            15'd14976: data <= 8'hFF;
            15'd14977: data <= 8'hFF;
            15'd14978: data <= 8'hFF;
            15'd14979: data <= 8'hF0;
            15'd14980: data <= 8'h7F;
            15'd14981: data <= 8'hFF;
            15'd14982: data <= 8'hFF;
            15'd14983: data <= 8'hFF;
            15'd14984: data <= 8'hFF;
            15'd14985: data <= 8'hFF;
            15'd14986: data <= 8'hFF;
            15'd14987: data <= 8'hFF;
            15'd14988: data <= 8'hFF;
            15'd14989: data <= 8'hFF;
            15'd14990: data <= 8'hFF;
            15'd14991: data <= 8'hFF;
            15'd14992: data <= 8'hFF;
            15'd14993: data <= 8'hF0;
            15'd14994: data <= 8'h00;
            15'd14995: data <= 8'h00;
            15'd14996: data <= 8'h00;
            15'd14997: data <= 8'h00;
            15'd14998: data <= 8'h00;
            15'd14999: data <= 8'h00;
            15'd15000: data <= 8'h00;
            15'd15001: data <= 8'h00;
            15'd15002: data <= 8'h00;
            15'd15003: data <= 8'h00;
            15'd15004: data <= 8'h00;
            15'd15005: data <= 8'h03;
            15'd15006: data <= 8'hFF;
            15'd15007: data <= 8'hFF;
            15'd15008: data <= 8'hFF;
            15'd15009: data <= 8'hF0;
            15'd15010: data <= 8'h7F;
            15'd15011: data <= 8'hFF;
            15'd15012: data <= 8'hFF;
            15'd15013: data <= 8'hFF;
            15'd15014: data <= 8'hFF;
            15'd15015: data <= 8'hFF;
            15'd15016: data <= 8'hFF;
            15'd15017: data <= 8'hFF;
            15'd15018: data <= 8'hFF;
            15'd15019: data <= 8'hFF;
            15'd15020: data <= 8'hFF;
            15'd15021: data <= 8'hFF;
            15'd15022: data <= 8'hFF;
            15'd15023: data <= 8'hF0;
            15'd15024: data <= 8'h00;
            15'd15025: data <= 8'h00;
            15'd15026: data <= 8'h00;
            15'd15027: data <= 8'h00;
            15'd15028: data <= 8'h00;
            15'd15029: data <= 8'h00;
            15'd15030: data <= 8'h00;
            15'd15031: data <= 8'h00;
            15'd15032: data <= 8'h00;
            15'd15033: data <= 8'h00;
            15'd15034: data <= 8'h00;
            15'd15035: data <= 8'h03;
            15'd15036: data <= 8'hFF;
            15'd15037: data <= 8'hFF;
            15'd15038: data <= 8'hFF;
            15'd15039: data <= 8'hF0;
            15'd15040: data <= 8'h7F;
            15'd15041: data <= 8'hFF;
            15'd15042: data <= 8'hFF;
            15'd15043: data <= 8'hFF;
            15'd15044: data <= 8'hFF;
            15'd15045: data <= 8'hFF;
            15'd15046: data <= 8'hFF;
            15'd15047: data <= 8'hFF;
            15'd15048: data <= 8'hFF;
            15'd15049: data <= 8'hFF;
            15'd15050: data <= 8'hFF;
            15'd15051: data <= 8'hFF;
            15'd15052: data <= 8'hFF;
            15'd15053: data <= 8'hF0;
            15'd15054: data <= 8'h00;
            15'd15055: data <= 8'h00;
            15'd15056: data <= 8'h00;
            15'd15057: data <= 8'h00;
            15'd15058: data <= 8'h00;
            15'd15059: data <= 8'h00;
            15'd15060: data <= 8'h00;
            15'd15061: data <= 8'h00;
            15'd15062: data <= 8'h00;
            15'd15063: data <= 8'h00;
            15'd15064: data <= 8'h00;
            15'd15065: data <= 8'h03;
            15'd15066: data <= 8'hFF;
            15'd15067: data <= 8'hFF;
            15'd15068: data <= 8'hFF;
            15'd15069: data <= 8'hF0;
            15'd15070: data <= 8'h7F;
            15'd15071: data <= 8'hFF;
            15'd15072: data <= 8'hFF;
            15'd15073: data <= 8'hFF;
            15'd15074: data <= 8'hFF;
            15'd15075: data <= 8'hFF;
            15'd15076: data <= 8'hFF;
            15'd15077: data <= 8'hFF;
            15'd15078: data <= 8'hFF;
            15'd15079: data <= 8'hFF;
            15'd15080: data <= 8'hFF;
            15'd15081: data <= 8'hFF;
            15'd15082: data <= 8'hFF;
            15'd15083: data <= 8'hF8;
            15'd15084: data <= 8'h00;
            15'd15085: data <= 8'h00;
            15'd15086: data <= 8'h00;
            15'd15087: data <= 8'h00;
            15'd15088: data <= 8'h00;
            15'd15089: data <= 8'h00;
            15'd15090: data <= 8'h00;
            15'd15091: data <= 8'h00;
            15'd15092: data <= 8'h00;
            15'd15093: data <= 8'h00;
            15'd15094: data <= 8'h00;
            15'd15095: data <= 8'h03;
            15'd15096: data <= 8'hFF;
            15'd15097: data <= 8'hFF;
            15'd15098: data <= 8'hFF;
            15'd15099: data <= 8'hE0;
            15'd15100: data <= 8'h7F;
            15'd15101: data <= 8'hFF;
            15'd15102: data <= 8'hFF;
            15'd15103: data <= 8'hFF;
            15'd15104: data <= 8'hFF;
            15'd15105: data <= 8'hFF;
            15'd15106: data <= 8'hFF;
            15'd15107: data <= 8'hFF;
            15'd15108: data <= 8'hFF;
            15'd15109: data <= 8'hFF;
            15'd15110: data <= 8'hFF;
            15'd15111: data <= 8'hFF;
            15'd15112: data <= 8'hFF;
            15'd15113: data <= 8'hF8;
            15'd15114: data <= 8'h00;
            15'd15115: data <= 8'h00;
            15'd15116: data <= 8'h00;
            15'd15117: data <= 8'h00;
            15'd15118: data <= 8'h00;
            15'd15119: data <= 8'h00;
            15'd15120: data <= 8'h00;
            15'd15121: data <= 8'h00;
            15'd15122: data <= 8'h00;
            15'd15123: data <= 8'h00;
            15'd15124: data <= 8'h00;
            15'd15125: data <= 8'h03;
            15'd15126: data <= 8'hFF;
            15'd15127: data <= 8'hFF;
            15'd15128: data <= 8'hFF;
            15'd15129: data <= 8'hE0;
            15'd15130: data <= 8'h7F;
            15'd15131: data <= 8'hFF;
            15'd15132: data <= 8'hFF;
            15'd15133: data <= 8'hFF;
            15'd15134: data <= 8'hFF;
            15'd15135: data <= 8'hFF;
            15'd15136: data <= 8'hFF;
            15'd15137: data <= 8'hFF;
            15'd15138: data <= 8'hFF;
            15'd15139: data <= 8'hFF;
            15'd15140: data <= 8'hFF;
            15'd15141: data <= 8'hFF;
            15'd15142: data <= 8'hFF;
            15'd15143: data <= 8'hF8;
            15'd15144: data <= 8'h00;
            15'd15145: data <= 8'h00;
            15'd15146: data <= 8'h00;
            15'd15147: data <= 8'h00;
            15'd15148: data <= 8'h00;
            15'd15149: data <= 8'h00;
            15'd15150: data <= 8'h00;
            15'd15151: data <= 8'h00;
            15'd15152: data <= 8'h00;
            15'd15153: data <= 8'h00;
            15'd15154: data <= 8'h00;
            15'd15155: data <= 8'h03;
            15'd15156: data <= 8'hFF;
            15'd15157: data <= 8'hFF;
            15'd15158: data <= 8'hFF;
            15'd15159: data <= 8'hE0;
            15'd15160: data <= 8'h7F;
            15'd15161: data <= 8'hFF;
            15'd15162: data <= 8'hFF;
            15'd15163: data <= 8'hFF;
            15'd15164: data <= 8'hFF;
            15'd15165: data <= 8'hFF;
            15'd15166: data <= 8'hFF;
            15'd15167: data <= 8'hFF;
            15'd15168: data <= 8'hFF;
            15'd15169: data <= 8'hFF;
            15'd15170: data <= 8'hFF;
            15'd15171: data <= 8'hFF;
            15'd15172: data <= 8'hFF;
            15'd15173: data <= 8'hF8;
            15'd15174: data <= 8'h00;
            15'd15175: data <= 8'h00;
            15'd15176: data <= 8'h00;
            15'd15177: data <= 8'h00;
            15'd15178: data <= 8'h00;
            15'd15179: data <= 8'h00;
            15'd15180: data <= 8'h00;
            15'd15181: data <= 8'h00;
            15'd15182: data <= 8'h00;
            15'd15183: data <= 8'h00;
            15'd15184: data <= 8'h00;
            15'd15185: data <= 8'h03;
            15'd15186: data <= 8'hFF;
            15'd15187: data <= 8'hFF;
            15'd15188: data <= 8'hFF;
            15'd15189: data <= 8'hE0;
            15'd15190: data <= 8'h7F;
            15'd15191: data <= 8'hFF;
            15'd15192: data <= 8'hFF;
            15'd15193: data <= 8'hFF;
            15'd15194: data <= 8'hFF;
            15'd15195: data <= 8'hFF;
            15'd15196: data <= 8'hFF;
            15'd15197: data <= 8'hFF;
            15'd15198: data <= 8'hFF;
            15'd15199: data <= 8'hFF;
            15'd15200: data <= 8'hFF;
            15'd15201: data <= 8'hFF;
            15'd15202: data <= 8'hFF;
            15'd15203: data <= 8'hF8;
            15'd15204: data <= 8'h00;
            15'd15205: data <= 8'h00;
            15'd15206: data <= 8'h00;
            15'd15207: data <= 8'h00;
            15'd15208: data <= 8'h00;
            15'd15209: data <= 8'h00;
            15'd15210: data <= 8'h00;
            15'd15211: data <= 8'h00;
            15'd15212: data <= 8'h00;
            15'd15213: data <= 8'h00;
            15'd15214: data <= 8'h00;
            15'd15215: data <= 8'h03;
            15'd15216: data <= 8'hFF;
            15'd15217: data <= 8'hFF;
            15'd15218: data <= 8'hFF;
            15'd15219: data <= 8'hF0;
            15'd15220: data <= 8'hFF;
            15'd15221: data <= 8'hFF;
            15'd15222: data <= 8'hFF;
            15'd15223: data <= 8'hFF;
            15'd15224: data <= 8'hFF;
            15'd15225: data <= 8'hFF;
            15'd15226: data <= 8'hFF;
            15'd15227: data <= 8'hFF;
            15'd15228: data <= 8'hFF;
            15'd15229: data <= 8'hFF;
            15'd15230: data <= 8'hFF;
            15'd15231: data <= 8'hFF;
            15'd15232: data <= 8'hFF;
            15'd15233: data <= 8'hFC;
            15'd15234: data <= 8'h00;
            15'd15235: data <= 8'h00;
            15'd15236: data <= 8'h00;
            15'd15237: data <= 8'h00;
            15'd15238: data <= 8'h00;
            15'd15239: data <= 8'h00;
            15'd15240: data <= 8'h00;
            15'd15241: data <= 8'h00;
            15'd15242: data <= 8'h00;
            15'd15243: data <= 8'h00;
            15'd15244: data <= 8'h00;
            15'd15245: data <= 8'h03;
            15'd15246: data <= 8'hFF;
            15'd15247: data <= 8'hFF;
            15'd15248: data <= 8'hFF;
            15'd15249: data <= 8'hFF;
            15'd15250: data <= 8'hFF;
            15'd15251: data <= 8'hFF;
            15'd15252: data <= 8'hFF;
            15'd15253: data <= 8'hFF;
            15'd15254: data <= 8'hFF;
            15'd15255: data <= 8'hFF;
            15'd15256: data <= 8'hFF;
            15'd15257: data <= 8'hFF;
            15'd15258: data <= 8'hFF;
            15'd15259: data <= 8'hFF;
            15'd15260: data <= 8'hFF;
            15'd15261: data <= 8'hFF;
            15'd15262: data <= 8'hFF;
            15'd15263: data <= 8'hFF;
            15'd15264: data <= 8'h80;
            15'd15265: data <= 8'h00;
            15'd15266: data <= 8'h00;
            15'd15267: data <= 8'h00;
            15'd15268: data <= 8'h00;
            15'd15269: data <= 8'h00;
            15'd15270: data <= 8'h00;
            15'd15271: data <= 8'h00;
            15'd15272: data <= 8'h00;
            15'd15273: data <= 8'h00;
            15'd15274: data <= 8'h00;
            15'd15275: data <= 8'h03;
            15'd15276: data <= 8'hFF;
            15'd15277: data <= 8'hFF;
            15'd15278: data <= 8'hFF;
            15'd15279: data <= 8'hFF;
            15'd15280: data <= 8'hFF;
            15'd15281: data <= 8'hFF;
            15'd15282: data <= 8'hFF;
            15'd15283: data <= 8'hFF;
            15'd15284: data <= 8'hFF;
            15'd15285: data <= 8'hFF;
            15'd15286: data <= 8'hFF;
            15'd15287: data <= 8'hFF;
            15'd15288: data <= 8'hFF;
            15'd15289: data <= 8'hFF;
            15'd15290: data <= 8'hFF;
            15'd15291: data <= 8'hFF;
            15'd15292: data <= 8'hFF;
            15'd15293: data <= 8'hFF;
            15'd15294: data <= 8'h80;
            15'd15295: data <= 8'h00;
            15'd15296: data <= 8'h00;
            15'd15297: data <= 8'h00;
            15'd15298: data <= 8'h00;
            15'd15299: data <= 8'h00;
            15'd15300: data <= 8'h00;
            15'd15301: data <= 8'h00;
            15'd15302: data <= 8'h00;
            15'd15303: data <= 8'h00;
            15'd15304: data <= 8'h00;
            15'd15305: data <= 8'h03;
            15'd15306: data <= 8'hFF;
            15'd15307: data <= 8'hFF;
            15'd15308: data <= 8'hFF;
            15'd15309: data <= 8'hFF;
            15'd15310: data <= 8'hFF;
            15'd15311: data <= 8'hFF;
            15'd15312: data <= 8'hFF;
            15'd15313: data <= 8'hFF;
            15'd15314: data <= 8'hFF;
            15'd15315: data <= 8'hFF;
            15'd15316: data <= 8'hFF;
            15'd15317: data <= 8'hFF;
            15'd15318: data <= 8'hFF;
            15'd15319: data <= 8'hFF;
            15'd15320: data <= 8'hFF;
            15'd15321: data <= 8'hFF;
            15'd15322: data <= 8'hFF;
            15'd15323: data <= 8'hFF;
            15'd15324: data <= 8'h80;
            15'd15325: data <= 8'h00;
            15'd15326: data <= 8'h00;
            15'd15327: data <= 8'h00;
            15'd15328: data <= 8'h00;
            15'd15329: data <= 8'h00;
            15'd15330: data <= 8'h00;
            15'd15331: data <= 8'h00;
            15'd15332: data <= 8'h00;
            15'd15333: data <= 8'h00;
            15'd15334: data <= 8'h00;
            15'd15335: data <= 8'h03;
            15'd15336: data <= 8'hFF;
            15'd15337: data <= 8'hFF;
            15'd15338: data <= 8'hFF;
            15'd15339: data <= 8'hFF;
            15'd15340: data <= 8'hFF;
            15'd15341: data <= 8'hFF;
            15'd15342: data <= 8'hFF;
            15'd15343: data <= 8'hFF;
            15'd15344: data <= 8'hFF;
            15'd15345: data <= 8'hFF;
            15'd15346: data <= 8'hFF;
            15'd15347: data <= 8'hFF;
            15'd15348: data <= 8'hFF;
            15'd15349: data <= 8'hFF;
            15'd15350: data <= 8'hFF;
            15'd15351: data <= 8'hFF;
            15'd15352: data <= 8'hFF;
            15'd15353: data <= 8'hFF;
            15'd15354: data <= 8'h80;
            15'd15355: data <= 8'h00;
            15'd15356: data <= 8'h00;
            15'd15357: data <= 8'h00;
            15'd15358: data <= 8'h00;
            15'd15359: data <= 8'h00;
            15'd15360: data <= 8'h00;
            15'd15361: data <= 8'h00;
            15'd15362: data <= 8'h00;
            15'd15363: data <= 8'h00;
            15'd15364: data <= 8'h00;
            15'd15365: data <= 8'h03;
            15'd15366: data <= 8'hFF;
            15'd15367: data <= 8'hFF;
            15'd15368: data <= 8'hFF;
            15'd15369: data <= 8'hFF;
            15'd15370: data <= 8'hFF;
            15'd15371: data <= 8'hFF;
            15'd15372: data <= 8'hFF;
            15'd15373: data <= 8'hFF;
            15'd15374: data <= 8'hFF;
            15'd15375: data <= 8'hFF;
            15'd15376: data <= 8'hFF;
            15'd15377: data <= 8'hFF;
            15'd15378: data <= 8'hFF;
            15'd15379: data <= 8'hFF;
            15'd15380: data <= 8'hFF;
            15'd15381: data <= 8'hFF;
            15'd15382: data <= 8'hFF;
            15'd15383: data <= 8'hFF;
            15'd15384: data <= 8'h80;
            15'd15385: data <= 8'h00;
            15'd15386: data <= 8'h00;
            15'd15387: data <= 8'h00;
            15'd15388: data <= 8'h00;
            15'd15389: data <= 8'h00;
            15'd15390: data <= 8'h00;
            15'd15391: data <= 8'h00;
            15'd15392: data <= 8'h00;
            15'd15393: data <= 8'h00;
            15'd15394: data <= 8'h00;
            15'd15395: data <= 8'h03;
            15'd15396: data <= 8'hFF;
            15'd15397: data <= 8'hFF;
            15'd15398: data <= 8'hFF;
            15'd15399: data <= 8'hFF;
            15'd15400: data <= 8'hFF;
            15'd15401: data <= 8'hFF;
            15'd15402: data <= 8'hFF;
            15'd15403: data <= 8'hFF;
            15'd15404: data <= 8'hFF;
            15'd15405: data <= 8'hFF;
            15'd15406: data <= 8'hFF;
            15'd15407: data <= 8'hFF;
            15'd15408: data <= 8'hFF;
            15'd15409: data <= 8'hFF;
            15'd15410: data <= 8'hFF;
            15'd15411: data <= 8'hFF;
            15'd15412: data <= 8'hFF;
            15'd15413: data <= 8'hFF;
            15'd15414: data <= 8'h80;
            15'd15415: data <= 8'h00;
            15'd15416: data <= 8'h00;
            15'd15417: data <= 8'h00;
            15'd15418: data <= 8'h00;
            15'd15419: data <= 8'h00;
            15'd15420: data <= 8'h00;
            15'd15421: data <= 8'h00;
            15'd15422: data <= 8'h00;
            15'd15423: data <= 8'h00;
            15'd15424: data <= 8'h00;
            15'd15425: data <= 8'h03;
            15'd15426: data <= 8'hFF;
            15'd15427: data <= 8'hFF;
            15'd15428: data <= 8'hFF;
            15'd15429: data <= 8'hFF;
            15'd15430: data <= 8'hFF;
            15'd15431: data <= 8'hFF;
            15'd15432: data <= 8'hFF;
            15'd15433: data <= 8'hFF;
            15'd15434: data <= 8'hFF;
            15'd15435: data <= 8'hFF;
            15'd15436: data <= 8'hFF;
            15'd15437: data <= 8'hFF;
            15'd15438: data <= 8'hFF;
            15'd15439: data <= 8'hFF;
            15'd15440: data <= 8'hFF;
            15'd15441: data <= 8'hFF;
            15'd15442: data <= 8'hFF;
            15'd15443: data <= 8'hFF;
            15'd15444: data <= 8'h80;
            15'd15445: data <= 8'h00;
            15'd15446: data <= 8'h00;
            15'd15447: data <= 8'h00;
            15'd15448: data <= 8'h00;
            15'd15449: data <= 8'h00;
            15'd15450: data <= 8'h00;
            15'd15451: data <= 8'h00;
            15'd15452: data <= 8'h00;
            15'd15453: data <= 8'h00;
            15'd15454: data <= 8'h00;
            15'd15455: data <= 8'h03;
            15'd15456: data <= 8'hFF;
            15'd15457: data <= 8'hFF;
            15'd15458: data <= 8'hFF;
            15'd15459: data <= 8'hFF;
            15'd15460: data <= 8'hFF;
            15'd15461: data <= 8'hFF;
            15'd15462: data <= 8'hFF;
            15'd15463: data <= 8'hFF;
            15'd15464: data <= 8'hFF;
            15'd15465: data <= 8'hFF;
            15'd15466: data <= 8'hFF;
            15'd15467: data <= 8'hFF;
            15'd15468: data <= 8'h8F;
            15'd15469: data <= 8'hFF;
            15'd15470: data <= 8'hFF;
            15'd15471: data <= 8'hFF;
            15'd15472: data <= 8'hFF;
            15'd15473: data <= 8'hFF;
            15'd15474: data <= 8'h80;
            15'd15475: data <= 8'h00;
            15'd15476: data <= 8'h00;
            15'd15477: data <= 8'h00;
            15'd15478: data <= 8'h00;
            15'd15479: data <= 8'h00;
            15'd15480: data <= 8'h00;
            15'd15481: data <= 8'h00;
            15'd15482: data <= 8'h00;
            15'd15483: data <= 8'h00;
            15'd15484: data <= 8'h00;
            15'd15485: data <= 8'h03;
            15'd15486: data <= 8'hFF;
            15'd15487: data <= 8'hFF;
            15'd15488: data <= 8'hFF;
            15'd15489: data <= 8'hFF;
            15'd15490: data <= 8'hFB;
            15'd15491: data <= 8'hFF;
            15'd15492: data <= 8'hFF;
            15'd15493: data <= 8'hFF;
            15'd15494: data <= 8'hFE;
            15'd15495: data <= 8'hFF;
            15'd15496: data <= 8'hFF;
            15'd15497: data <= 8'hF8;
            15'd15498: data <= 8'h07;
            15'd15499: data <= 8'hFF;
            15'd15500: data <= 8'hFF;
            15'd15501: data <= 8'hFF;
            15'd15502: data <= 8'hFF;
            15'd15503: data <= 8'hFF;
            15'd15504: data <= 8'h80;
            15'd15505: data <= 8'h00;
            15'd15506: data <= 8'h00;
            15'd15507: data <= 8'h00;
            15'd15508: data <= 8'h00;
            15'd15509: data <= 8'h00;
            15'd15510: data <= 8'h00;
            15'd15511: data <= 8'h00;
            15'd15512: data <= 8'h00;
            15'd15513: data <= 8'h00;
            15'd15514: data <= 8'h00;
            15'd15515: data <= 8'h03;
            15'd15516: data <= 8'hFF;
            15'd15517: data <= 8'hE0;
            15'd15518: data <= 8'h00;
            15'd15519: data <= 8'h3C;
            15'd15520: data <= 8'h0B;
            15'd15521: data <= 8'h7F;
            15'd15522: data <= 8'hFF;
            15'd15523: data <= 8'hFF;
            15'd15524: data <= 8'hFC;
            15'd15525: data <= 8'h7F;
            15'd15526: data <= 8'hFF;
            15'd15527: data <= 8'hC3;
            15'd15528: data <= 8'hF1;
            15'd15529: data <= 8'hFF;
            15'd15530: data <= 8'hFF;
            15'd15531: data <= 8'hE0;
            15'd15532: data <= 8'h1F;
            15'd15533: data <= 8'hFF;
            15'd15534: data <= 8'h80;
            15'd15535: data <= 8'h00;
            15'd15536: data <= 8'h00;
            15'd15537: data <= 8'h00;
            15'd15538: data <= 8'h00;
            15'd15539: data <= 8'h00;
            15'd15540: data <= 8'h00;
            15'd15541: data <= 8'h00;
            15'd15542: data <= 8'h00;
            15'd15543: data <= 8'h00;
            15'd15544: data <= 8'h00;
            15'd15545: data <= 8'h03;
            15'd15546: data <= 8'hFF;
            15'd15547: data <= 8'hFF;
            15'd15548: data <= 8'h77;
            15'd15549: data <= 8'hF0;
            15'd15550: data <= 8'h7B;
            15'd15551: data <= 8'h1F;
            15'd15552: data <= 8'hFF;
            15'd15553: data <= 8'hFE;
            15'd15554: data <= 8'h00;
            15'd15555: data <= 8'h00;
            15'd15556: data <= 8'hFF;
            15'd15557: data <= 8'h9F;
            15'd15558: data <= 8'hFC;
            15'd15559: data <= 8'h3F;
            15'd15560: data <= 8'hF8;
            15'd15561: data <= 8'h7F;
            15'd15562: data <= 8'h9F;
            15'd15563: data <= 8'hFF;
            15'd15564: data <= 8'h80;
            15'd15565: data <= 8'h00;
            15'd15566: data <= 8'h00;
            15'd15567: data <= 8'h00;
            15'd15568: data <= 8'h00;
            15'd15569: data <= 8'h00;
            15'd15570: data <= 8'h00;
            15'd15571: data <= 8'h00;
            15'd15572: data <= 8'h00;
            15'd15573: data <= 8'h00;
            15'd15574: data <= 8'h00;
            15'd15575: data <= 8'h03;
            15'd15576: data <= 8'hFF;
            15'd15577: data <= 8'hFF;
            15'd15578: data <= 8'h77;
            15'd15579: data <= 8'hFE;
            15'd15580: data <= 8'h7B;
            15'd15581: data <= 8'hDF;
            15'd15582: data <= 8'hFF;
            15'd15583: data <= 8'hFF;
            15'd15584: data <= 8'hFE;
            15'd15585: data <= 8'hFF;
            15'd15586: data <= 8'hFF;
            15'd15587: data <= 8'h3F;
            15'd15588: data <= 8'hFF;
            15'd15589: data <= 8'h9F;
            15'd15590: data <= 8'hFB;
            15'd15591: data <= 8'h37;
            15'd15592: data <= 8'h9F;
            15'd15593: data <= 8'hFF;
            15'd15594: data <= 8'h80;
            15'd15595: data <= 8'h00;
            15'd15596: data <= 8'h00;
            15'd15597: data <= 8'h00;
            15'd15598: data <= 8'h00;
            15'd15599: data <= 8'h00;
            15'd15600: data <= 8'h00;
            15'd15601: data <= 8'h00;
            15'd15602: data <= 8'h00;
            15'd15603: data <= 8'h00;
            15'd15604: data <= 8'h00;
            15'd15605: data <= 8'h03;
            15'd15606: data <= 8'hFF;
            15'd15607: data <= 8'hF0;
            15'd15608: data <= 8'h00;
            15'd15609: data <= 8'h3E;
            15'd15610: data <= 8'h7B;
            15'd15611: data <= 8'hFF;
            15'd15612: data <= 8'hFF;
            15'd15613: data <= 8'hFF;
            15'd15614: data <= 8'hC0;
            15'd15615: data <= 8'h0F;
            15'd15616: data <= 8'hFE;
            15'd15617: data <= 8'h7F;
            15'd15618: data <= 8'hFF;
            15'd15619: data <= 8'h9F;
            15'd15620: data <= 8'hFB;
            15'd15621: data <= 8'h37;
            15'd15622: data <= 8'h9F;
            15'd15623: data <= 8'hFF;
            15'd15624: data <= 8'h80;
            15'd15625: data <= 8'h00;
            15'd15626: data <= 8'h00;
            15'd15627: data <= 8'h00;
            15'd15628: data <= 8'h00;
            15'd15629: data <= 8'h00;
            15'd15630: data <= 8'h00;
            15'd15631: data <= 8'h00;
            15'd15632: data <= 8'h00;
            15'd15633: data <= 8'h00;
            15'd15634: data <= 8'h00;
            15'd15635: data <= 8'h03;
            15'd15636: data <= 8'hFF;
            15'd15637: data <= 8'hE7;
            15'd15638: data <= 8'h77;
            15'd15639: data <= 8'h30;
            15'd15640: data <= 8'h00;
            15'd15641: data <= 8'h0F;
            15'd15642: data <= 8'hFF;
            15'd15643: data <= 8'hFF;
            15'd15644: data <= 8'h80;
            15'd15645: data <= 8'h03;
            15'd15646: data <= 8'hFE;
            15'd15647: data <= 8'hEF;
            15'd15648: data <= 8'hFF;
            15'd15649: data <= 8'hDF;
            15'd15650: data <= 8'hFB;
            15'd15651: data <= 8'h27;
            15'd15652: data <= 8'h9F;
            15'd15653: data <= 8'hFF;
            15'd15654: data <= 8'h80;
            15'd15655: data <= 8'h00;
            15'd15656: data <= 8'h00;
            15'd15657: data <= 8'h00;
            15'd15658: data <= 8'h00;
            15'd15659: data <= 8'h00;
            15'd15660: data <= 8'h00;
            15'd15661: data <= 8'h00;
            15'd15662: data <= 8'h00;
            15'd15663: data <= 8'h00;
            15'd15664: data <= 8'h00;
            15'd15665: data <= 8'h03;
            15'd15666: data <= 8'hFF;
            15'd15667: data <= 8'hE7;
            15'd15668: data <= 8'h77;
            15'd15669: data <= 8'h30;
            15'd15670: data <= 8'h00;
            15'd15671: data <= 8'h07;
            15'd15672: data <= 8'hFF;
            15'd15673: data <= 8'hFF;
            15'd15674: data <= 8'h9F;
            15'd15675: data <= 8'hF3;
            15'd15676: data <= 8'hFE;
            15'd15677: data <= 8'hFF;
            15'd15678: data <= 8'hFF;
            15'd15679: data <= 8'hCF;
            15'd15680: data <= 8'hFB;
            15'd15681: data <= 8'h27;
            15'd15682: data <= 8'hBF;
            15'd15683: data <= 8'hFF;
            15'd15684: data <= 8'h80;
            15'd15685: data <= 8'h00;
            15'd15686: data <= 8'h00;
            15'd15687: data <= 8'h00;
            15'd15688: data <= 8'h00;
            15'd15689: data <= 8'h00;
            15'd15690: data <= 8'h00;
            15'd15691: data <= 8'h00;
            15'd15692: data <= 8'h00;
            15'd15693: data <= 8'h00;
            15'd15694: data <= 8'h00;
            15'd15695: data <= 8'h03;
            15'd15696: data <= 8'hFF;
            15'd15697: data <= 8'hE0;
            15'd15698: data <= 8'h00;
            15'd15699: data <= 8'h3E;
            15'd15700: data <= 8'h79;
            15'd15701: data <= 8'hFC;
            15'd15702: data <= 8'h00;
            15'd15703: data <= 8'h03;
            15'd15704: data <= 8'h80;
            15'd15705: data <= 8'h03;
            15'd15706: data <= 8'hFE;
            15'd15707: data <= 8'hFF;
            15'd15708: data <= 8'hFF;
            15'd15709: data <= 8'hE7;
            15'd15710: data <= 8'hFB;
            15'd15711: data <= 8'h27;
            15'd15712: data <= 8'hBF;
            15'd15713: data <= 8'hFF;
            15'd15714: data <= 8'h80;
            15'd15715: data <= 8'h00;
            15'd15716: data <= 8'h00;
            15'd15717: data <= 8'h00;
            15'd15718: data <= 8'h00;
            15'd15719: data <= 8'h00;
            15'd15720: data <= 8'h00;
            15'd15721: data <= 8'h00;
            15'd15722: data <= 8'h00;
            15'd15723: data <= 8'h00;
            15'd15724: data <= 8'h00;
            15'd15725: data <= 8'h03;
            15'd15726: data <= 8'hFF;
            15'd15727: data <= 8'hF7;
            15'd15728: data <= 8'h7F;
            15'd15729: data <= 8'h3E;
            15'd15730: data <= 8'h79;
            15'd15731: data <= 8'hC8;
            15'd15732: data <= 8'h00;
            15'd15733: data <= 8'h03;
            15'd15734: data <= 8'h9F;
            15'd15735: data <= 8'hF3;
            15'd15736: data <= 8'hFE;
            15'd15737: data <= 8'hE3;
            15'd15738: data <= 8'hFF;
            15'd15739: data <= 8'hF7;
            15'd15740: data <= 8'hFB;
            15'd15741: data <= 8'h20;
            15'd15742: data <= 8'h0F;
            15'd15743: data <= 8'hFF;
            15'd15744: data <= 8'h80;
            15'd15745: data <= 8'h00;
            15'd15746: data <= 8'h00;
            15'd15747: data <= 8'h00;
            15'd15748: data <= 8'h00;
            15'd15749: data <= 8'h00;
            15'd15750: data <= 8'h00;
            15'd15751: data <= 8'h00;
            15'd15752: data <= 8'h00;
            15'd15753: data <= 8'h00;
            15'd15754: data <= 8'h00;
            15'd15755: data <= 8'h03;
            15'd15756: data <= 8'hFF;
            15'd15757: data <= 8'hFF;
            15'd15758: data <= 8'h7F;
            15'd15759: data <= 8'hFE;
            15'd15760: data <= 8'h0D;
            15'd15761: data <= 8'h9F;
            15'd15762: data <= 8'hFF;
            15'd15763: data <= 8'hFF;
            15'd15764: data <= 8'h9F;
            15'd15765: data <= 8'hF3;
            15'd15766: data <= 8'hFE;
            15'd15767: data <= 8'h05;
            15'd15768: data <= 8'hFF;
            15'd15769: data <= 8'hF3;
            15'd15770: data <= 8'hFB;
            15'd15771: data <= 8'h3F;
            15'd15772: data <= 8'hEF;
            15'd15773: data <= 8'hFF;
            15'd15774: data <= 8'h80;
            15'd15775: data <= 8'h00;
            15'd15776: data <= 8'h00;
            15'd15777: data <= 8'h00;
            15'd15778: data <= 8'h00;
            15'd15779: data <= 8'h00;
            15'd15780: data <= 8'h00;
            15'd15781: data <= 8'h00;
            15'd15782: data <= 8'h00;
            15'd15783: data <= 8'h00;
            15'd15784: data <= 8'h00;
            15'd15785: data <= 8'h03;
            15'd15786: data <= 8'hFF;
            15'd15787: data <= 8'hC0;
            15'd15788: data <= 8'h00;
            15'd15789: data <= 8'h10;
            15'd15790: data <= 8'h1D;
            15'd15791: data <= 8'h3F;
            15'd15792: data <= 8'hFF;
            15'd15793: data <= 8'hFF;
            15'd15794: data <= 8'h80;
            15'd15795: data <= 8'h03;
            15'd15796: data <= 8'hFF;
            15'd15797: data <= 8'h01;
            15'd15798: data <= 8'hFF;
            15'd15799: data <= 8'hFB;
            15'd15800: data <= 8'hFB;
            15'd15801: data <= 8'h3F;
            15'd15802: data <= 8'hEF;
            15'd15803: data <= 8'hFF;
            15'd15804: data <= 8'h80;
            15'd15805: data <= 8'h00;
            15'd15806: data <= 8'h00;
            15'd15807: data <= 8'h00;
            15'd15808: data <= 8'h00;
            15'd15809: data <= 8'h00;
            15'd15810: data <= 8'h00;
            15'd15811: data <= 8'h00;
            15'd15812: data <= 8'h00;
            15'd15813: data <= 8'h00;
            15'd15814: data <= 8'h00;
            15'd15815: data <= 8'h03;
            15'd15816: data <= 8'hFF;
            15'd15817: data <= 8'hFC;
            15'd15818: data <= 8'hF9;
            15'd15819: data <= 8'hF2;
            15'd15820: data <= 8'h7C;
            15'd15821: data <= 8'h7F;
            15'd15822: data <= 8'hFF;
            15'd15823: data <= 8'hFF;
            15'd15824: data <= 8'h9F;
            15'd15825: data <= 8'hF3;
            15'd15826: data <= 8'hFF;
            15'd15827: data <= 8'h9F;
            15'd15828: data <= 8'hFF;
            15'd15829: data <= 8'hFB;
            15'd15830: data <= 8'hFB;
            15'd15831: data <= 8'h3F;
            15'd15832: data <= 8'hEF;
            15'd15833: data <= 8'hFF;
            15'd15834: data <= 8'h80;
            15'd15835: data <= 8'h00;
            15'd15836: data <= 8'h00;
            15'd15837: data <= 8'h00;
            15'd15838: data <= 8'h00;
            15'd15839: data <= 8'h00;
            15'd15840: data <= 8'h00;
            15'd15841: data <= 8'h00;
            15'd15842: data <= 8'h00;
            15'd15843: data <= 8'h00;
            15'd15844: data <= 8'h00;
            15'd15845: data <= 8'h03;
            15'd15846: data <= 8'hFF;
            15'd15847: data <= 8'hFD;
            15'd15848: data <= 8'hFB;
            15'd15849: data <= 8'hFE;
            15'd15850: data <= 8'h7C;
            15'd15851: data <= 8'hFF;
            15'd15852: data <= 8'hFF;
            15'd15853: data <= 8'hFF;
            15'd15854: data <= 8'h80;
            15'd15855: data <= 8'h03;
            15'd15856: data <= 8'hFF;
            15'd15857: data <= 8'hAD;
            15'd15858: data <= 8'hFF;
            15'd15859: data <= 8'hF9;
            15'd15860: data <= 8'hF8;
            15'd15861: data <= 8'h00;
            15'd15862: data <= 8'h2F;
            15'd15863: data <= 8'hFF;
            15'd15864: data <= 8'h80;
            15'd15865: data <= 8'h00;
            15'd15866: data <= 8'h00;
            15'd15867: data <= 8'h00;
            15'd15868: data <= 8'h00;
            15'd15869: data <= 8'h00;
            15'd15870: data <= 8'h00;
            15'd15871: data <= 8'h00;
            15'd15872: data <= 8'h00;
            15'd15873: data <= 8'h00;
            15'd15874: data <= 8'h00;
            15'd15875: data <= 8'h03;
            15'd15876: data <= 8'hFF;
            15'd15877: data <= 8'hFC;
            15'd15878: data <= 8'h27;
            15'd15879: data <= 8'hFE;
            15'd15880: data <= 8'h70;
            15'd15881: data <= 8'hE7;
            15'd15882: data <= 8'hFF;
            15'd15883: data <= 8'hFF;
            15'd15884: data <= 8'h80;
            15'd15885: data <= 8'h03;
            15'd15886: data <= 8'hFF;
            15'd15887: data <= 8'hAE;
            15'd15888: data <= 8'h67;
            15'd15889: data <= 8'hFD;
            15'd15890: data <= 8'hFB;
            15'd15891: data <= 8'h3F;
            15'd15892: data <= 8'hEF;
            15'd15893: data <= 8'hFF;
            15'd15894: data <= 8'h80;
            15'd15895: data <= 8'h00;
            15'd15896: data <= 8'h00;
            15'd15897: data <= 8'h00;
            15'd15898: data <= 8'h00;
            15'd15899: data <= 8'h00;
            15'd15900: data <= 8'h00;
            15'd15901: data <= 8'h00;
            15'd15902: data <= 8'h00;
            15'd15903: data <= 8'h00;
            15'd15904: data <= 8'h00;
            15'd15905: data <= 8'h03;
            15'd15906: data <= 8'hFF;
            15'd15907: data <= 8'hFF;
            15'd15908: data <= 8'h87;
            15'd15909: data <= 8'hFE;
            15'd15910: data <= 8'h66;
            15'd15911: data <= 8'h6F;
            15'd15912: data <= 8'hFF;
            15'd15913: data <= 8'hFF;
            15'd15914: data <= 8'h9F;
            15'd15915: data <= 8'hF3;
            15'd15916: data <= 8'hFF;
            15'd15917: data <= 8'hB7;
            15'd15918: data <= 8'h8F;
            15'd15919: data <= 8'hFC;
            15'd15920: data <= 8'hFF;
            15'd15921: data <= 8'hFF;
            15'd15922: data <= 8'hEF;
            15'd15923: data <= 8'hFF;
            15'd15924: data <= 8'h80;
            15'd15925: data <= 8'h00;
            15'd15926: data <= 8'h00;
            15'd15927: data <= 8'h00;
            15'd15928: data <= 8'h00;
            15'd15929: data <= 8'h00;
            15'd15930: data <= 8'h00;
            15'd15931: data <= 8'h00;
            15'd15932: data <= 8'h00;
            15'd15933: data <= 8'h00;
            15'd15934: data <= 8'h00;
            15'd15935: data <= 8'h03;
            15'd15936: data <= 8'hFF;
            15'd15937: data <= 8'hFC;
            15'd15938: data <= 8'h30;
            15'd15939: data <= 8'h7E;
            15'd15940: data <= 8'h4F;
            15'd15941: data <= 8'h2F;
            15'd15942: data <= 8'hFF;
            15'd15943: data <= 8'hFE;
            15'd15944: data <= 8'h00;
            15'd15945: data <= 8'h00;
            15'd15946: data <= 8'hFF;
            15'd15947: data <= 8'hF7;
            15'd15948: data <= 8'hFF;
            15'd15949: data <= 8'hFC;
            15'd15950: data <= 8'hFF;
            15'd15951: data <= 8'hFC;
            15'd15952: data <= 8'h0F;
            15'd15953: data <= 8'hFF;
            15'd15954: data <= 8'h80;
            15'd15955: data <= 8'h00;
            15'd15956: data <= 8'h00;
            15'd15957: data <= 8'h00;
            15'd15958: data <= 8'h00;
            15'd15959: data <= 8'h00;
            15'd15960: data <= 8'h00;
            15'd15961: data <= 8'h00;
            15'd15962: data <= 8'h00;
            15'd15963: data <= 8'h00;
            15'd15964: data <= 8'h00;
            15'd15965: data <= 8'h03;
            15'd15966: data <= 8'hFF;
            15'd15967: data <= 8'hE1;
            15'd15968: data <= 8'hFE;
            15'd15969: data <= 8'h38;
            15'd15970: data <= 8'hFF;
            15'd15971: data <= 8'h8F;
            15'd15972: data <= 8'hFF;
            15'd15973: data <= 8'hFE;
            15'd15974: data <= 8'h00;
            15'd15975: data <= 8'h00;
            15'd15976: data <= 8'hFF;
            15'd15977: data <= 8'hFB;
            15'd15978: data <= 8'hFF;
            15'd15979: data <= 8'hFE;
            15'd15980: data <= 8'hFF;
            15'd15981: data <= 8'hFC;
            15'd15982: data <= 8'h1F;
            15'd15983: data <= 8'hFF;
            15'd15984: data <= 8'h80;
            15'd15985: data <= 8'h00;
            15'd15986: data <= 8'h00;
            15'd15987: data <= 8'h00;
            15'd15988: data <= 8'h00;
            15'd15989: data <= 8'h00;
            15'd15990: data <= 8'h00;
            15'd15991: data <= 8'h00;
            15'd15992: data <= 8'h00;
            15'd15993: data <= 8'h00;
            15'd15994: data <= 8'h00;
            15'd15995: data <= 8'h03;
            15'd15996: data <= 8'hFF;
            15'd15997: data <= 8'hFF;
            15'd15998: data <= 8'hFF;
            15'd15999: data <= 8'hFF;
            15'd16000: data <= 8'hFF;
            15'd16001: data <= 8'hFF;
            15'd16002: data <= 8'hFF;
            15'd16003: data <= 8'hFF;
            15'd16004: data <= 8'hFF;
            15'd16005: data <= 8'hFF;
            15'd16006: data <= 8'hFF;
            15'd16007: data <= 8'hBD;
            15'd16008: data <= 8'hFF;
            15'd16009: data <= 8'hFE;
            15'd16010: data <= 8'hFF;
            15'd16011: data <= 8'hFF;
            15'd16012: data <= 8'hFF;
            15'd16013: data <= 8'hFF;
            15'd16014: data <= 8'h80;
            15'd16015: data <= 8'h00;
            15'd16016: data <= 8'h00;
            15'd16017: data <= 8'h00;
            15'd16018: data <= 8'h00;
            15'd16019: data <= 8'h00;
            15'd16020: data <= 8'h00;
            15'd16021: data <= 8'h00;
            15'd16022: data <= 8'h00;
            15'd16023: data <= 8'h00;
            15'd16024: data <= 8'h00;
            15'd16025: data <= 8'h03;
            15'd16026: data <= 8'hFF;
            15'd16027: data <= 8'hFF;
            15'd16028: data <= 8'hFF;
            15'd16029: data <= 8'hFF;
            15'd16030: data <= 8'hFF;
            15'd16031: data <= 8'hFF;
            15'd16032: data <= 8'hFF;
            15'd16033: data <= 8'hFF;
            15'd16034: data <= 8'hFF;
            15'd16035: data <= 8'hFF;
            15'd16036: data <= 8'hFF;
            15'd16037: data <= 8'hBE;
            15'd16038: data <= 8'h7F;
            15'd16039: data <= 8'hFE;
            15'd16040: data <= 8'h7F;
            15'd16041: data <= 8'hFF;
            15'd16042: data <= 8'hFF;
            15'd16043: data <= 8'hFF;
            15'd16044: data <= 8'h80;
            15'd16045: data <= 8'h00;
            15'd16046: data <= 8'h00;
            15'd16047: data <= 8'h00;
            15'd16048: data <= 8'h00;
            15'd16049: data <= 8'h00;
            15'd16050: data <= 8'h00;
            15'd16051: data <= 8'h00;
            15'd16052: data <= 8'h00;
            15'd16053: data <= 8'h00;
            15'd16054: data <= 8'h00;
            15'd16055: data <= 8'h03;
            15'd16056: data <= 8'hFF;
            15'd16057: data <= 8'hFF;
            15'd16058: data <= 8'hFF;
            15'd16059: data <= 8'hFF;
            15'd16060: data <= 8'hFF;
            15'd16061: data <= 8'hFF;
            15'd16062: data <= 8'hFF;
            15'd16063: data <= 8'hFF;
            15'd16064: data <= 8'hFF;
            15'd16065: data <= 8'hFF;
            15'd16066: data <= 8'hFF;
            15'd16067: data <= 8'hBF;
            15'd16068: data <= 8'h03;
            15'd16069: data <= 8'hFE;
            15'd16070: data <= 8'h7F;
            15'd16071: data <= 8'hFF;
            15'd16072: data <= 8'hFF;
            15'd16073: data <= 8'hFF;
            15'd16074: data <= 8'h80;
            15'd16075: data <= 8'h00;
            15'd16076: data <= 8'h00;
            15'd16077: data <= 8'h00;
            15'd16078: data <= 8'h00;
            15'd16079: data <= 8'h00;
            15'd16080: data <= 8'h00;
            15'd16081: data <= 8'h00;
            15'd16082: data <= 8'h00;
            15'd16083: data <= 8'h00;
            15'd16084: data <= 8'h00;
            15'd16085: data <= 8'h03;
            15'd16086: data <= 8'hFF;
            15'd16087: data <= 8'hFF;
            15'd16088: data <= 8'hFF;
            15'd16089: data <= 8'hFF;
            15'd16090: data <= 8'hFF;
            15'd16091: data <= 8'hFF;
            15'd16092: data <= 8'hFF;
            15'd16093: data <= 8'hFF;
            15'd16094: data <= 8'hFF;
            15'd16095: data <= 8'hFF;
            15'd16096: data <= 8'hFF;
            15'd16097: data <= 8'hBF;
            15'd16098: data <= 8'hFF;
            15'd16099: data <= 8'hFF;
            15'd16100: data <= 8'h7F;
            15'd16101: data <= 8'hFF;
            15'd16102: data <= 8'hFF;
            15'd16103: data <= 8'hFF;
            15'd16104: data <= 8'h80;
            15'd16105: data <= 8'h00;
            15'd16106: data <= 8'h00;
            15'd16107: data <= 8'h00;
            15'd16108: data <= 8'h00;
            15'd16109: data <= 8'h00;
            15'd16110: data <= 8'h00;
            15'd16111: data <= 8'h00;
            15'd16112: data <= 8'h00;
            15'd16113: data <= 8'h00;
            15'd16114: data <= 8'h00;
            15'd16115: data <= 8'h03;
            15'd16116: data <= 8'hFF;
            15'd16117: data <= 8'hFF;
            15'd16118: data <= 8'hFF;
            15'd16119: data <= 8'hFF;
            15'd16120: data <= 8'hFF;
            15'd16121: data <= 8'hFF;
            15'd16122: data <= 8'hFF;
            15'd16123: data <= 8'hFF;
            15'd16124: data <= 8'hFF;
            15'd16125: data <= 8'hFF;
            15'd16126: data <= 8'hFF;
            15'd16127: data <= 8'hBF;
            15'd16128: data <= 8'hFF;
            15'd16129: data <= 8'hFF;
            15'd16130: data <= 8'h7F;
            15'd16131: data <= 8'hFF;
            15'd16132: data <= 8'hFF;
            15'd16133: data <= 8'hFF;
            15'd16134: data <= 8'h80;
            15'd16135: data <= 8'h00;
            15'd16136: data <= 8'h00;
            15'd16137: data <= 8'h00;
            15'd16138: data <= 8'h00;
            15'd16139: data <= 8'h00;
            15'd16140: data <= 8'h00;
            15'd16141: data <= 8'h00;
            15'd16142: data <= 8'h00;
            15'd16143: data <= 8'h00;
            15'd16144: data <= 8'h00;
            15'd16145: data <= 8'h03;
            15'd16146: data <= 8'hFF;
            15'd16147: data <= 8'hFF;
            15'd16148: data <= 8'hFF;
            15'd16149: data <= 8'hFF;
            15'd16150: data <= 8'hFF;
            15'd16151: data <= 8'hFF;
            15'd16152: data <= 8'hFF;
            15'd16153: data <= 8'hFF;
            15'd16154: data <= 8'hFF;
            15'd16155: data <= 8'hFF;
            15'd16156: data <= 8'hFF;
            15'd16157: data <= 8'hBF;
            15'd16158: data <= 8'hFF;
            15'd16159: data <= 8'hFF;
            15'd16160: data <= 8'hFF;
            15'd16161: data <= 8'hFF;
            15'd16162: data <= 8'hFF;
            15'd16163: data <= 8'hFF;
            15'd16164: data <= 8'h80;
            15'd16165: data <= 8'h00;
            15'd16166: data <= 8'h00;
            15'd16167: data <= 8'h00;
            15'd16168: data <= 8'h00;
            15'd16169: data <= 8'h00;
            15'd16170: data <= 8'h00;
            15'd16171: data <= 8'h00;
            15'd16172: data <= 8'h00;
            15'd16173: data <= 8'h00;
            15'd16174: data <= 8'h00;
            15'd16175: data <= 8'h03;
            15'd16176: data <= 8'hFF;
            15'd16177: data <= 8'hFF;
            15'd16178: data <= 8'hFF;
            15'd16179: data <= 8'hFF;
            15'd16180: data <= 8'hFF;
            15'd16181: data <= 8'hFF;
            15'd16182: data <= 8'hFF;
            15'd16183: data <= 8'hFF;
            15'd16184: data <= 8'hFF;
            15'd16185: data <= 8'hFF;
            15'd16186: data <= 8'hFF;
            15'd16187: data <= 8'hFF;
            15'd16188: data <= 8'hFF;
            15'd16189: data <= 8'hFF;
            15'd16190: data <= 8'hFF;
            15'd16191: data <= 8'hFF;
            15'd16192: data <= 8'hFF;
            15'd16193: data <= 8'hFF;
            15'd16194: data <= 8'h80;
            15'd16195: data <= 8'h00;
            15'd16196: data <= 8'h00;
            15'd16197: data <= 8'h00;
            15'd16198: data <= 8'h00;
            15'd16199: data <= 8'h00;
            15'd16200: data <= 8'h00;
            15'd16201: data <= 8'h00;
            15'd16202: data <= 8'h00;
            15'd16203: data <= 8'h00;
            15'd16204: data <= 8'h00;
            15'd16205: data <= 8'h03;
            15'd16206: data <= 8'hFF;
            15'd16207: data <= 8'hFF;
            15'd16208: data <= 8'hFF;
            15'd16209: data <= 8'hFF;
            15'd16210: data <= 8'hFF;
            15'd16211: data <= 8'hFF;
            15'd16212: data <= 8'hFF;
            15'd16213: data <= 8'hFF;
            15'd16214: data <= 8'hFF;
            15'd16215: data <= 8'hFF;
            15'd16216: data <= 8'hFF;
            15'd16217: data <= 8'hFF;
            15'd16218: data <= 8'hFF;
            15'd16219: data <= 8'hFF;
            15'd16220: data <= 8'hFF;
            15'd16221: data <= 8'hFF;
            15'd16222: data <= 8'hFF;
            15'd16223: data <= 8'hFF;
            15'd16224: data <= 8'h80;
            15'd16225: data <= 8'h00;
            15'd16226: data <= 8'h00;
            15'd16227: data <= 8'h00;
            15'd16228: data <= 8'h00;
            15'd16229: data <= 8'h00;
            15'd16230: data <= 8'h00;
            15'd16231: data <= 8'h00;
            15'd16232: data <= 8'h00;
            15'd16233: data <= 8'h00;
            15'd16234: data <= 8'h00;
            15'd16235: data <= 8'h03;
            15'd16236: data <= 8'hFF;
            15'd16237: data <= 8'hFF;
            15'd16238: data <= 8'hFF;
            15'd16239: data <= 8'hFF;
            15'd16240: data <= 8'hFF;
            15'd16241: data <= 8'hFF;
            15'd16242: data <= 8'hFF;
            15'd16243: data <= 8'hFF;
            15'd16244: data <= 8'hFF;
            15'd16245: data <= 8'hFF;
            15'd16246: data <= 8'hFF;
            15'd16247: data <= 8'hFF;
            15'd16248: data <= 8'hFF;
            15'd16249: data <= 8'hFF;
            15'd16250: data <= 8'hFF;
            15'd16251: data <= 8'hFF;
            15'd16252: data <= 8'hFF;
            15'd16253: data <= 8'hFF;
            15'd16254: data <= 8'h80;
            15'd16255: data <= 8'h00;
            15'd16256: data <= 8'h00;
            15'd16257: data <= 8'h00;
            15'd16258: data <= 8'h00;
            15'd16259: data <= 8'h00;
            15'd16260: data <= 8'h00;
            15'd16261: data <= 8'h00;
            15'd16262: data <= 8'h00;
            15'd16263: data <= 8'h00;
            15'd16264: data <= 8'h00;
            15'd16265: data <= 8'h03;
            15'd16266: data <= 8'hFF;
            15'd16267: data <= 8'hFF;
            15'd16268: data <= 8'hFF;
            15'd16269: data <= 8'hFF;
            15'd16270: data <= 8'hFF;
            15'd16271: data <= 8'hFF;
            15'd16272: data <= 8'hFF;
            15'd16273: data <= 8'hFF;
            15'd16274: data <= 8'hFF;
            15'd16275: data <= 8'hFF;
            15'd16276: data <= 8'hFF;
            15'd16277: data <= 8'hFF;
            15'd16278: data <= 8'hFF;
            15'd16279: data <= 8'hFF;
            15'd16280: data <= 8'hFF;
            15'd16281: data <= 8'hFF;
            15'd16282: data <= 8'hFF;
            15'd16283: data <= 8'hFF;
            15'd16284: data <= 8'h80;
            15'd16285: data <= 8'h00;
            15'd16286: data <= 8'h00;
            15'd16287: data <= 8'h00;
            15'd16288: data <= 8'h00;
            15'd16289: data <= 8'h00;
            15'd16290: data <= 8'h00;
            15'd16291: data <= 8'h00;
            15'd16292: data <= 8'h00;
            15'd16293: data <= 8'h00;
            15'd16294: data <= 8'h00;
            15'd16295: data <= 8'h03;
            15'd16296: data <= 8'hFF;
            15'd16297: data <= 8'hFF;
            15'd16298: data <= 8'hFF;
            15'd16299: data <= 8'hFF;
            15'd16300: data <= 8'hFF;
            15'd16301: data <= 8'hFF;
            15'd16302: data <= 8'hFF;
            15'd16303: data <= 8'hFF;
            15'd16304: data <= 8'hFF;
            15'd16305: data <= 8'hFF;
            15'd16306: data <= 8'hFF;
            15'd16307: data <= 8'hFF;
            15'd16308: data <= 8'hFF;
            15'd16309: data <= 8'hFF;
            15'd16310: data <= 8'hFF;
            15'd16311: data <= 8'hFF;
            15'd16312: data <= 8'hFF;
            15'd16313: data <= 8'hFF;
            15'd16314: data <= 8'h80;
            15'd16315: data <= 8'h00;
            15'd16316: data <= 8'h00;
            15'd16317: data <= 8'h00;
            15'd16318: data <= 8'h00;
            15'd16319: data <= 8'h00;
            15'd16320: data <= 8'h00;
            15'd16321: data <= 8'h00;
            15'd16322: data <= 8'h00;
            15'd16323: data <= 8'h00;
            15'd16324: data <= 8'h00;
            15'd16325: data <= 8'h03;
            15'd16326: data <= 8'hFF;
            15'd16327: data <= 8'hFF;
            15'd16328: data <= 8'hFF;
            15'd16329: data <= 8'hFF;
            15'd16330: data <= 8'hFF;
            15'd16331: data <= 8'hFF;
            15'd16332: data <= 8'hFF;
            15'd16333: data <= 8'hFF;
            15'd16334: data <= 8'hFF;
            15'd16335: data <= 8'hFF;
            15'd16336: data <= 8'hFF;
            15'd16337: data <= 8'hFF;
            15'd16338: data <= 8'hFF;
            15'd16339: data <= 8'hFF;
            15'd16340: data <= 8'hFF;
            15'd16341: data <= 8'hFF;
            15'd16342: data <= 8'hFF;
            15'd16343: data <= 8'hFF;
            15'd16344: data <= 8'h80;
            15'd16345: data <= 8'h00;
            15'd16346: data <= 8'h00;
            15'd16347: data <= 8'h00;
            15'd16348: data <= 8'h00;
            15'd16349: data <= 8'h00;
            15'd16350: data <= 8'h00;
            15'd16351: data <= 8'h00;
            15'd16352: data <= 8'h00;
            15'd16353: data <= 8'h00;
            15'd16354: data <= 8'h00;
            15'd16355: data <= 8'h03;
            15'd16356: data <= 8'hFF;
            15'd16357: data <= 8'hFF;
            15'd16358: data <= 8'hFF;
            15'd16359: data <= 8'hFF;
            15'd16360: data <= 8'hFF;
            15'd16361: data <= 8'hFF;
            15'd16362: data <= 8'hFF;
            15'd16363: data <= 8'hFF;
            15'd16364: data <= 8'hFF;
            15'd16365: data <= 8'hFF;
            15'd16366: data <= 8'hFF;
            15'd16367: data <= 8'hFF;
            15'd16368: data <= 8'hFF;
            15'd16369: data <= 8'hFF;
            15'd16370: data <= 8'hFF;
            15'd16371: data <= 8'hFF;
            15'd16372: data <= 8'hFF;
            15'd16373: data <= 8'hFF;
            15'd16374: data <= 8'h80;
            15'd16375: data <= 8'h00;
            15'd16376: data <= 8'h00;
            15'd16377: data <= 8'h00;
            15'd16378: data <= 8'h00;
            15'd16379: data <= 8'h00;
            15'd16380: data <= 8'h00;
            15'd16381: data <= 8'h00;
            15'd16382: data <= 8'h00;
            15'd16383: data <= 8'h00;
            15'd16384: data <= 8'h00;
            15'd16385: data <= 8'h03;
            15'd16386: data <= 8'hFF;
            15'd16387: data <= 8'hFF;
            15'd16388: data <= 8'hFF;
            15'd16389: data <= 8'hFF;
            15'd16390: data <= 8'hFF;
            15'd16391: data <= 8'hFF;
            15'd16392: data <= 8'hFF;
            15'd16393: data <= 8'hFF;
            15'd16394: data <= 8'hFF;
            15'd16395: data <= 8'hFF;
            15'd16396: data <= 8'hFF;
            15'd16397: data <= 8'hFF;
            15'd16398: data <= 8'hFF;
            15'd16399: data <= 8'hFF;
            15'd16400: data <= 8'hFF;
            15'd16401: data <= 8'hFF;
            15'd16402: data <= 8'hFF;
            15'd16403: data <= 8'hFF;
            15'd16404: data <= 8'h80;
            15'd16405: data <= 8'h00;
            15'd16406: data <= 8'h00;
            15'd16407: data <= 8'h00;
            15'd16408: data <= 8'h00;
            15'd16409: data <= 8'h00;
            15'd16410: data <= 8'h00;
            15'd16411: data <= 8'h00;
            15'd16412: data <= 8'h00;
            15'd16413: data <= 8'h00;
            15'd16414: data <= 8'h00;
            15'd16415: data <= 8'h03;
            15'd16416: data <= 8'hFF;
            15'd16417: data <= 8'hFF;
            15'd16418: data <= 8'hFF;
            15'd16419: data <= 8'hFF;
            15'd16420: data <= 8'hFF;
            15'd16421: data <= 8'hFF;
            15'd16422: data <= 8'hFF;
            15'd16423: data <= 8'hFF;
            15'd16424: data <= 8'hFF;
            15'd16425: data <= 8'hFF;
            15'd16426: data <= 8'hFF;
            15'd16427: data <= 8'hFF;
            15'd16428: data <= 8'hFF;
            15'd16429: data <= 8'hFF;
            15'd16430: data <= 8'hFF;
            15'd16431: data <= 8'hFF;
            15'd16432: data <= 8'hFF;
            15'd16433: data <= 8'hFF;
            15'd16434: data <= 8'h80;
            15'd16435: data <= 8'h00;
            15'd16436: data <= 8'h00;
            15'd16437: data <= 8'h00;
            15'd16438: data <= 8'h00;
            15'd16439: data <= 8'h00;
            15'd16440: data <= 8'h00;
            15'd16441: data <= 8'h00;
            15'd16442: data <= 8'h00;
            15'd16443: data <= 8'h00;
            15'd16444: data <= 8'h00;
            15'd16445: data <= 8'h03;
            15'd16446: data <= 8'hFF;
            15'd16447: data <= 8'hFF;
            15'd16448: data <= 8'hFF;
            15'd16449: data <= 8'hFF;
            15'd16450: data <= 8'hFF;
            15'd16451: data <= 8'hFF;
            15'd16452: data <= 8'hFF;
            15'd16453: data <= 8'hFF;
            15'd16454: data <= 8'hFF;
            15'd16455: data <= 8'hFF;
            15'd16456: data <= 8'hFF;
            15'd16457: data <= 8'hFF;
            15'd16458: data <= 8'hFF;
            15'd16459: data <= 8'hFF;
            15'd16460: data <= 8'hFF;
            15'd16461: data <= 8'hFF;
            15'd16462: data <= 8'hFF;
            15'd16463: data <= 8'hFF;
            15'd16464: data <= 8'h80;
            15'd16465: data <= 8'h00;
            15'd16466: data <= 8'h00;
            15'd16467: data <= 8'h00;
            15'd16468: data <= 8'h00;
            15'd16469: data <= 8'h00;
            15'd16470: data <= 8'h00;
            15'd16471: data <= 8'h00;
            15'd16472: data <= 8'h00;
            15'd16473: data <= 8'h00;
            15'd16474: data <= 8'h00;
            15'd16475: data <= 8'h03;
            15'd16476: data <= 8'hFF;
            15'd16477: data <= 8'hFF;
            15'd16478: data <= 8'hFF;
            15'd16479: data <= 8'hFF;
            15'd16480: data <= 8'hFF;
            15'd16481: data <= 8'hFF;
            15'd16482: data <= 8'hFF;
            15'd16483: data <= 8'hFF;
            15'd16484: data <= 8'hFF;
            15'd16485: data <= 8'hFF;
            15'd16486: data <= 8'hFF;
            15'd16487: data <= 8'hFF;
            15'd16488: data <= 8'hFF;
            15'd16489: data <= 8'hFF;
            15'd16490: data <= 8'hFF;
            15'd16491: data <= 8'hFF;
            15'd16492: data <= 8'hFF;
            15'd16493: data <= 8'hFF;
            15'd16494: data <= 8'h80;
            15'd16495: data <= 8'h00;
            15'd16496: data <= 8'h00;
            15'd16497: data <= 8'h00;
            15'd16498: data <= 8'h00;
            15'd16499: data <= 8'h00;
            15'd16500: data <= 8'h00;
            15'd16501: data <= 8'h00;
            15'd16502: data <= 8'h00;
            15'd16503: data <= 8'h00;
            15'd16504: data <= 8'h00;
            15'd16505: data <= 8'h03;
            15'd16506: data <= 8'hFF;
            15'd16507: data <= 8'hFF;
            15'd16508: data <= 8'hFF;
            15'd16509: data <= 8'hFF;
            15'd16510: data <= 8'hFF;
            15'd16511: data <= 8'hFF;
            15'd16512: data <= 8'hFF;
            15'd16513: data <= 8'hFF;
            15'd16514: data <= 8'hFF;
            15'd16515: data <= 8'hFF;
            15'd16516: data <= 8'hFF;
            15'd16517: data <= 8'hFF;
            15'd16518: data <= 8'hFF;
            15'd16519: data <= 8'hFF;
            15'd16520: data <= 8'hFF;
            15'd16521: data <= 8'hFF;
            15'd16522: data <= 8'hFF;
            15'd16523: data <= 8'hFF;
            15'd16524: data <= 8'h80;
            15'd16525: data <= 8'h00;
            15'd16526: data <= 8'h00;
            15'd16527: data <= 8'h00;
            15'd16528: data <= 8'h00;
            15'd16529: data <= 8'h00;
            15'd16530: data <= 8'h00;
            15'd16531: data <= 8'h00;
            15'd16532: data <= 8'h00;
            15'd16533: data <= 8'h00;
            15'd16534: data <= 8'h00;
            15'd16535: data <= 8'h03;
            15'd16536: data <= 8'hFF;
            15'd16537: data <= 8'hFF;
            15'd16538: data <= 8'hFF;
            15'd16539: data <= 8'hFF;
            15'd16540: data <= 8'hFF;
            15'd16541: data <= 8'hFF;
            15'd16542: data <= 8'hFF;
            15'd16543: data <= 8'hFF;
            15'd16544: data <= 8'hFF;
            15'd16545: data <= 8'hFF;
            15'd16546: data <= 8'hFF;
            15'd16547: data <= 8'hFF;
            15'd16548: data <= 8'hFF;
            15'd16549: data <= 8'hFF;
            15'd16550: data <= 8'hFF;
            15'd16551: data <= 8'hFF;
            15'd16552: data <= 8'hFF;
            15'd16553: data <= 8'hFF;
            15'd16554: data <= 8'h80;
            15'd16555: data <= 8'h00;
            15'd16556: data <= 8'h00;
            15'd16557: data <= 8'h00;
            15'd16558: data <= 8'h00;
            15'd16559: data <= 8'h00;
            15'd16560: data <= 8'h00;
            15'd16561: data <= 8'h00;
            15'd16562: data <= 8'h00;
            15'd16563: data <= 8'h00;
            15'd16564: data <= 8'h00;
            15'd16565: data <= 8'h03;
            15'd16566: data <= 8'hFF;
            15'd16567: data <= 8'hFF;
            15'd16568: data <= 8'hFF;
            15'd16569: data <= 8'hFF;
            15'd16570: data <= 8'hFF;
            15'd16571: data <= 8'hFF;
            15'd16572: data <= 8'hFF;
            15'd16573: data <= 8'hFF;
            15'd16574: data <= 8'hFF;
            15'd16575: data <= 8'hFF;
            15'd16576: data <= 8'hFF;
            15'd16577: data <= 8'hFF;
            15'd16578: data <= 8'hFF;
            15'd16579: data <= 8'hFF;
            15'd16580: data <= 8'hFF;
            15'd16581: data <= 8'hFF;
            15'd16582: data <= 8'hFF;
            15'd16583: data <= 8'hFF;
            15'd16584: data <= 8'h80;
            15'd16585: data <= 8'h00;
            15'd16586: data <= 8'h00;
            15'd16587: data <= 8'h00;
            15'd16588: data <= 8'h00;
            15'd16589: data <= 8'h00;
            15'd16590: data <= 8'h00;
            15'd16591: data <= 8'h00;
            15'd16592: data <= 8'h00;
            15'd16593: data <= 8'h00;
            15'd16594: data <= 8'h00;
            15'd16595: data <= 8'h03;
            15'd16596: data <= 8'hFF;
            15'd16597: data <= 8'hFF;
            15'd16598: data <= 8'hFF;
            15'd16599: data <= 8'hFF;
            15'd16600: data <= 8'hFF;
            15'd16601: data <= 8'hFF;
            15'd16602: data <= 8'hFF;
            15'd16603: data <= 8'hFF;
            15'd16604: data <= 8'hFF;
            15'd16605: data <= 8'hFF;
            15'd16606: data <= 8'hFF;
            15'd16607: data <= 8'hFF;
            15'd16608: data <= 8'hFF;
            15'd16609: data <= 8'hFF;
            15'd16610: data <= 8'hFF;
            15'd16611: data <= 8'hFF;
            15'd16612: data <= 8'hFF;
            15'd16613: data <= 8'hFF;
            15'd16614: data <= 8'h80;
            15'd16615: data <= 8'h00;
            15'd16616: data <= 8'h00;
            15'd16617: data <= 8'h00;
            15'd16618: data <= 8'h00;
            15'd16619: data <= 8'h00;
            15'd16620: data <= 8'h00;
            15'd16621: data <= 8'h00;
            15'd16622: data <= 8'h00;
            15'd16623: data <= 8'h00;
            15'd16624: data <= 8'h00;
            15'd16625: data <= 8'h03;
            15'd16626: data <= 8'hFF;
            15'd16627: data <= 8'hFF;
            15'd16628: data <= 8'hFF;
            15'd16629: data <= 8'hFF;
            15'd16630: data <= 8'hFF;
            15'd16631: data <= 8'hFF;
            15'd16632: data <= 8'hFF;
            15'd16633: data <= 8'hFF;
            15'd16634: data <= 8'hFF;
            15'd16635: data <= 8'hFF;
            15'd16636: data <= 8'hFF;
            15'd16637: data <= 8'hFF;
            15'd16638: data <= 8'hFF;
            15'd16639: data <= 8'hFF;
            15'd16640: data <= 8'hFF;
            15'd16641: data <= 8'hFF;
            15'd16642: data <= 8'hFF;
            15'd16643: data <= 8'hFF;
            15'd16644: data <= 8'h80;
            15'd16645: data <= 8'h00;
            15'd16646: data <= 8'h00;
            15'd16647: data <= 8'h00;
            15'd16648: data <= 8'h00;
            15'd16649: data <= 8'h00;
            15'd16650: data <= 8'h00;
            15'd16651: data <= 8'h00;
            15'd16652: data <= 8'h00;
            15'd16653: data <= 8'h00;
            15'd16654: data <= 8'h00;
            15'd16655: data <= 8'h03;
            15'd16656: data <= 8'hFF;
            15'd16657: data <= 8'hFF;
            15'd16658: data <= 8'hFF;
            15'd16659: data <= 8'hFF;
            15'd16660: data <= 8'hFF;
            15'd16661: data <= 8'hFF;
            15'd16662: data <= 8'hFF;
            15'd16663: data <= 8'hFF;
            15'd16664: data <= 8'hFF;
            15'd16665: data <= 8'hFF;
            15'd16666: data <= 8'hFF;
            15'd16667: data <= 8'hFF;
            15'd16668: data <= 8'hFF;
            15'd16669: data <= 8'hFF;
            15'd16670: data <= 8'hFF;
            15'd16671: data <= 8'hFF;
            15'd16672: data <= 8'hFF;
            15'd16673: data <= 8'hFF;
            15'd16674: data <= 8'h80;
            15'd16675: data <= 8'h00;
            15'd16676: data <= 8'h00;
            15'd16677: data <= 8'h00;
            15'd16678: data <= 8'h00;
            15'd16679: data <= 8'h00;
            15'd16680: data <= 8'h00;
            15'd16681: data <= 8'h00;
            15'd16682: data <= 8'h00;
            15'd16683: data <= 8'h00;
            15'd16684: data <= 8'h00;
            15'd16685: data <= 8'h03;
            15'd16686: data <= 8'hFF;
            15'd16687: data <= 8'hFF;
            15'd16688: data <= 8'hFF;
            15'd16689: data <= 8'hFF;
            15'd16690: data <= 8'hFF;
            15'd16691: data <= 8'hFF;
            15'd16692: data <= 8'hFF;
            15'd16693: data <= 8'hFF;
            15'd16694: data <= 8'hFF;
            15'd16695: data <= 8'hFF;
            15'd16696: data <= 8'hFF;
            15'd16697: data <= 8'hFF;
            15'd16698: data <= 8'hFF;
            15'd16699: data <= 8'hFF;
            15'd16700: data <= 8'hFF;
            15'd16701: data <= 8'hFF;
            15'd16702: data <= 8'hFF;
            15'd16703: data <= 8'hFF;
            15'd16704: data <= 8'h80;
            15'd16705: data <= 8'h00;
            15'd16706: data <= 8'h00;
            15'd16707: data <= 8'h00;
            15'd16708: data <= 8'h00;
            15'd16709: data <= 8'h00;
            15'd16710: data <= 8'h00;
            15'd16711: data <= 8'h00;
            15'd16712: data <= 8'h00;
            15'd16713: data <= 8'h00;
            15'd16714: data <= 8'h00;
            15'd16715: data <= 8'h03;
            15'd16716: data <= 8'hFF;
            15'd16717: data <= 8'hFF;
            15'd16718: data <= 8'hFF;
            15'd16719: data <= 8'hFF;
            15'd16720: data <= 8'hFF;
            15'd16721: data <= 8'hFF;
            15'd16722: data <= 8'hFF;
            15'd16723: data <= 8'hFF;
            15'd16724: data <= 8'hFF;
            15'd16725: data <= 8'hFF;
            15'd16726: data <= 8'hFF;
            15'd16727: data <= 8'hFF;
            15'd16728: data <= 8'hFF;
            15'd16729: data <= 8'hFF;
            15'd16730: data <= 8'hFF;
            15'd16731: data <= 8'hFF;
            15'd16732: data <= 8'hFF;
            15'd16733: data <= 8'hFF;
            15'd16734: data <= 8'h80;
            15'd16735: data <= 8'h00;
            15'd16736: data <= 8'h00;
            15'd16737: data <= 8'h00;
            15'd16738: data <= 8'h00;
            15'd16739: data <= 8'h00;
            15'd16740: data <= 8'h00;
            15'd16741: data <= 8'h00;
            15'd16742: data <= 8'h00;
            15'd16743: data <= 8'h00;
            15'd16744: data <= 8'h00;
            15'd16745: data <= 8'h03;
            15'd16746: data <= 8'hFF;
            15'd16747: data <= 8'hFF;
            15'd16748: data <= 8'hFF;
            15'd16749: data <= 8'hFF;
            15'd16750: data <= 8'hFF;
            15'd16751: data <= 8'hFF;
            15'd16752: data <= 8'hFF;
            15'd16753: data <= 8'hFF;
            15'd16754: data <= 8'hFF;
            15'd16755: data <= 8'hFF;
            15'd16756: data <= 8'hFF;
            15'd16757: data <= 8'hFF;
            15'd16758: data <= 8'hFF;
            15'd16759: data <= 8'hFF;
            15'd16760: data <= 8'hFF;
            15'd16761: data <= 8'hFF;
            15'd16762: data <= 8'hFF;
            15'd16763: data <= 8'hFF;
            15'd16764: data <= 8'h80;
            15'd16765: data <= 8'h00;
            15'd16766: data <= 8'h00;
            15'd16767: data <= 8'h00;
            15'd16768: data <= 8'h00;
            15'd16769: data <= 8'h00;
            15'd16770: data <= 8'h00;
            15'd16771: data <= 8'h00;
            15'd16772: data <= 8'h00;
            15'd16773: data <= 8'h00;
            15'd16774: data <= 8'h00;
            15'd16775: data <= 8'h03;
            15'd16776: data <= 8'hFF;
            15'd16777: data <= 8'hFF;
            15'd16778: data <= 8'hFF;
            15'd16779: data <= 8'hFF;
            15'd16780: data <= 8'hFF;
            15'd16781: data <= 8'hFF;
            15'd16782: data <= 8'hFF;
            15'd16783: data <= 8'hFF;
            15'd16784: data <= 8'hFF;
            15'd16785: data <= 8'hFF;
            15'd16786: data <= 8'hFF;
            15'd16787: data <= 8'hFF;
            15'd16788: data <= 8'hFF;
            15'd16789: data <= 8'hFF;
            15'd16790: data <= 8'hFF;
            15'd16791: data <= 8'hFF;
            15'd16792: data <= 8'hFF;
            15'd16793: data <= 8'hFF;
            15'd16794: data <= 8'h80;
            15'd16795: data <= 8'h00;
            15'd16796: data <= 8'h00;
            15'd16797: data <= 8'h00;
            15'd16798: data <= 8'h00;
            15'd16799: data <= 8'h00;
            15'd16800: data <= 8'h00;
            15'd16801: data <= 8'h00;
            15'd16802: data <= 8'h00;
            15'd16803: data <= 8'h00;
            15'd16804: data <= 8'h00;
            15'd16805: data <= 8'h03;
            15'd16806: data <= 8'hFF;
            15'd16807: data <= 8'hFF;
            15'd16808: data <= 8'hFF;
            15'd16809: data <= 8'hFF;
            15'd16810: data <= 8'hFF;
            15'd16811: data <= 8'hFF;
            15'd16812: data <= 8'hFF;
            15'd16813: data <= 8'hFF;
            15'd16814: data <= 8'hFF;
            15'd16815: data <= 8'hFF;
            15'd16816: data <= 8'hFF;
            15'd16817: data <= 8'hFF;
            15'd16818: data <= 8'hFF;
            15'd16819: data <= 8'hFF;
            15'd16820: data <= 8'hFF;
            15'd16821: data <= 8'hFF;
            15'd16822: data <= 8'hFF;
            15'd16823: data <= 8'hFF;
            15'd16824: data <= 8'h80;
            15'd16825: data <= 8'h00;
            15'd16826: data <= 8'h00;
            15'd16827: data <= 8'h00;
            15'd16828: data <= 8'h00;
            15'd16829: data <= 8'h00;
            15'd16830: data <= 8'h00;
            15'd16831: data <= 8'h00;
            15'd16832: data <= 8'h00;
            15'd16833: data <= 8'h00;
            15'd16834: data <= 8'h00;
            15'd16835: data <= 8'h03;
            15'd16836: data <= 8'hFF;
            15'd16837: data <= 8'hFF;
            15'd16838: data <= 8'hFF;
            15'd16839: data <= 8'hFF;
            15'd16840: data <= 8'hFF;
            15'd16841: data <= 8'hFF;
            15'd16842: data <= 8'hFF;
            15'd16843: data <= 8'hFF;
            15'd16844: data <= 8'hFF;
            15'd16845: data <= 8'hFF;
            15'd16846: data <= 8'hFF;
            15'd16847: data <= 8'hFF;
            15'd16848: data <= 8'hFF;
            15'd16849: data <= 8'hFF;
            15'd16850: data <= 8'hFF;
            15'd16851: data <= 8'hFF;
            15'd16852: data <= 8'hFF;
            15'd16853: data <= 8'hFF;
            15'd16854: data <= 8'h80;
            15'd16855: data <= 8'h00;
            15'd16856: data <= 8'h00;
            15'd16857: data <= 8'h00;
            15'd16858: data <= 8'h00;
            15'd16859: data <= 8'h00;
            15'd16860: data <= 8'h00;
            15'd16861: data <= 8'h00;
            15'd16862: data <= 8'h00;
            15'd16863: data <= 8'h00;
            15'd16864: data <= 8'h00;
            15'd16865: data <= 8'h03;
            15'd16866: data <= 8'hFF;
            15'd16867: data <= 8'hFF;
            15'd16868: data <= 8'hFF;
            15'd16869: data <= 8'hFF;
            15'd16870: data <= 8'hFF;
            15'd16871: data <= 8'hFF;
            15'd16872: data <= 8'hFF;
            15'd16873: data <= 8'hFF;
            15'd16874: data <= 8'hFF;
            15'd16875: data <= 8'hFF;
            15'd16876: data <= 8'hFF;
            15'd16877: data <= 8'hFF;
            15'd16878: data <= 8'hFF;
            15'd16879: data <= 8'hFF;
            15'd16880: data <= 8'hFF;
            15'd16881: data <= 8'hFF;
            15'd16882: data <= 8'hFF;
            15'd16883: data <= 8'hFF;
            15'd16884: data <= 8'h80;
            15'd16885: data <= 8'h00;
            15'd16886: data <= 8'h00;
            15'd16887: data <= 8'h00;
            15'd16888: data <= 8'h00;
            15'd16889: data <= 8'h00;
            15'd16890: data <= 8'h00;
            15'd16891: data <= 8'h00;
            15'd16892: data <= 8'h00;
            15'd16893: data <= 8'h00;
            15'd16894: data <= 8'h00;
            15'd16895: data <= 8'h03;
            15'd16896: data <= 8'hFF;
            15'd16897: data <= 8'hFF;
            15'd16898: data <= 8'hFF;
            15'd16899: data <= 8'hFF;
            15'd16900: data <= 8'hFF;
            15'd16901: data <= 8'hFF;
            15'd16902: data <= 8'hFF;
            15'd16903: data <= 8'hFF;
            15'd16904: data <= 8'hFF;
            15'd16905: data <= 8'hFF;
            15'd16906: data <= 8'hFF;
            15'd16907: data <= 8'hFF;
            15'd16908: data <= 8'hFF;
            15'd16909: data <= 8'hFF;
            15'd16910: data <= 8'hFF;
            15'd16911: data <= 8'hFF;
            15'd16912: data <= 8'hFF;
            15'd16913: data <= 8'hFF;
            15'd16914: data <= 8'h80;
            15'd16915: data <= 8'h00;
            15'd16916: data <= 8'h00;
            15'd16917: data <= 8'h00;
            15'd16918: data <= 8'h00;
            15'd16919: data <= 8'h00;
            15'd16920: data <= 8'h00;
            15'd16921: data <= 8'h00;
            15'd16922: data <= 8'h00;
            15'd16923: data <= 8'h00;
            15'd16924: data <= 8'h00;
            15'd16925: data <= 8'h03;
            15'd16926: data <= 8'hFF;
            15'd16927: data <= 8'hFF;
            15'd16928: data <= 8'hFF;
            15'd16929: data <= 8'hFF;
            15'd16930: data <= 8'hFF;
            15'd16931: data <= 8'hFF;
            15'd16932: data <= 8'hFF;
            15'd16933: data <= 8'hFF;
            15'd16934: data <= 8'hFF;
            15'd16935: data <= 8'hFF;
            15'd16936: data <= 8'hFF;
            15'd16937: data <= 8'hFF;
            15'd16938: data <= 8'hFF;
            15'd16939: data <= 8'hFF;
            15'd16940: data <= 8'hFF;
            15'd16941: data <= 8'hFF;
            15'd16942: data <= 8'hFF;
            15'd16943: data <= 8'hFF;
            15'd16944: data <= 8'h80;
            15'd16945: data <= 8'h00;
            15'd16946: data <= 8'h00;
            15'd16947: data <= 8'h00;
            15'd16948: data <= 8'h00;
            15'd16949: data <= 8'h00;
            15'd16950: data <= 8'h00;
            15'd16951: data <= 8'h00;
            15'd16952: data <= 8'h00;
            15'd16953: data <= 8'h00;
            15'd16954: data <= 8'h00;
            15'd16955: data <= 8'h03;
            15'd16956: data <= 8'hFF;
            15'd16957: data <= 8'hFF;
            15'd16958: data <= 8'hFF;
            15'd16959: data <= 8'hFF;
            15'd16960: data <= 8'hFF;
            15'd16961: data <= 8'hFF;
            15'd16962: data <= 8'hFF;
            15'd16963: data <= 8'hFF;
            15'd16964: data <= 8'hFF;
            15'd16965: data <= 8'hFF;
            15'd16966: data <= 8'hFF;
            15'd16967: data <= 8'hFF;
            15'd16968: data <= 8'hFF;
            15'd16969: data <= 8'hFF;
            15'd16970: data <= 8'hFF;
            15'd16971: data <= 8'hFF;
            15'd16972: data <= 8'hFF;
            15'd16973: data <= 8'hFF;
            15'd16974: data <= 8'h80;
            15'd16975: data <= 8'h00;
            15'd16976: data <= 8'h00;
            15'd16977: data <= 8'h00;
            15'd16978: data <= 8'h00;
            15'd16979: data <= 8'h00;
            15'd16980: data <= 8'h00;
            15'd16981: data <= 8'h00;
            15'd16982: data <= 8'h00;
            15'd16983: data <= 8'h00;
            15'd16984: data <= 8'h00;
            15'd16985: data <= 8'h03;
            15'd16986: data <= 8'hFF;
            15'd16987: data <= 8'hFF;
            15'd16988: data <= 8'hFF;
            15'd16989: data <= 8'hFF;
            15'd16990: data <= 8'hFF;
            15'd16991: data <= 8'hFF;
            15'd16992: data <= 8'hFF;
            15'd16993: data <= 8'hFF;
            15'd16994: data <= 8'hFF;
            15'd16995: data <= 8'hFF;
            15'd16996: data <= 8'hFF;
            15'd16997: data <= 8'hFF;
            15'd16998: data <= 8'hFF;
            15'd16999: data <= 8'hFF;
            15'd17000: data <= 8'hFF;
            15'd17001: data <= 8'hFF;
            15'd17002: data <= 8'hFF;
            15'd17003: data <= 8'hFF;
            15'd17004: data <= 8'h80;
            15'd17005: data <= 8'h00;
            15'd17006: data <= 8'h00;
            15'd17007: data <= 8'h00;
            15'd17008: data <= 8'h00;
            15'd17009: data <= 8'h00;
            15'd17010: data <= 8'h00;
            15'd17011: data <= 8'h00;
            15'd17012: data <= 8'h00;
            15'd17013: data <= 8'h00;
            15'd17014: data <= 8'h00;
            15'd17015: data <= 8'h03;
            15'd17016: data <= 8'hFF;
            15'd17017: data <= 8'hFF;
            15'd17018: data <= 8'hFF;
            15'd17019: data <= 8'hFF;
            15'd17020: data <= 8'hFF;
            15'd17021: data <= 8'hFF;
            15'd17022: data <= 8'hFF;
            15'd17023: data <= 8'hFF;
            15'd17024: data <= 8'hFF;
            15'd17025: data <= 8'hFF;
            15'd17026: data <= 8'hFF;
            15'd17027: data <= 8'hFF;
            15'd17028: data <= 8'hFF;
            15'd17029: data <= 8'hFF;
            15'd17030: data <= 8'hFF;
            15'd17031: data <= 8'hFF;
            15'd17032: data <= 8'hFF;
            15'd17033: data <= 8'hFF;
            15'd17034: data <= 8'h80;
            15'd17035: data <= 8'h00;
            15'd17036: data <= 8'h00;
            15'd17037: data <= 8'h00;
            15'd17038: data <= 8'h00;
            15'd17039: data <= 8'h00;
            15'd17040: data <= 8'h00;
            15'd17041: data <= 8'h00;
            15'd17042: data <= 8'h00;
            15'd17043: data <= 8'h00;
            15'd17044: data <= 8'h00;
            15'd17045: data <= 8'h03;
            15'd17046: data <= 8'hFF;
            15'd17047: data <= 8'hFF;
            15'd17048: data <= 8'hFF;
            15'd17049: data <= 8'hFF;
            15'd17050: data <= 8'hFF;
            15'd17051: data <= 8'hFF;
            15'd17052: data <= 8'hFF;
            15'd17053: data <= 8'hFF;
            15'd17054: data <= 8'hFF;
            15'd17055: data <= 8'hFF;
            15'd17056: data <= 8'hFF;
            15'd17057: data <= 8'hFF;
            15'd17058: data <= 8'hFF;
            15'd17059: data <= 8'hFF;
            15'd17060: data <= 8'hFF;
            15'd17061: data <= 8'hFF;
            15'd17062: data <= 8'hFF;
            15'd17063: data <= 8'hFF;
            15'd17064: data <= 8'h80;
            15'd17065: data <= 8'h00;
            15'd17066: data <= 8'h00;
            15'd17067: data <= 8'h00;
            15'd17068: data <= 8'h00;
            15'd17069: data <= 8'h00;
            15'd17070: data <= 8'h00;
            15'd17071: data <= 8'h00;
            15'd17072: data <= 8'h00;
            15'd17073: data <= 8'h00;
            15'd17074: data <= 8'h00;
            15'd17075: data <= 8'h03;
            15'd17076: data <= 8'hFF;
            15'd17077: data <= 8'hFF;
            15'd17078: data <= 8'hFF;
            15'd17079: data <= 8'hFF;
            15'd17080: data <= 8'hFF;
            15'd17081: data <= 8'hFF;
            15'd17082: data <= 8'hFF;
            15'd17083: data <= 8'hFF;
            15'd17084: data <= 8'hFF;
            15'd17085: data <= 8'hFF;
            15'd17086: data <= 8'hFF;
            15'd17087: data <= 8'hFF;
            15'd17088: data <= 8'hFF;
            15'd17089: data <= 8'hFF;
            15'd17090: data <= 8'hFF;
            15'd17091: data <= 8'hFF;
            15'd17092: data <= 8'hFF;
            15'd17093: data <= 8'hFF;
            15'd17094: data <= 8'h80;
            15'd17095: data <= 8'h00;
            15'd17096: data <= 8'h00;
            15'd17097: data <= 8'h00;
            15'd17098: data <= 8'h00;
            15'd17099: data <= 8'h00;
            15'd17100: data <= 8'h00;
            15'd17101: data <= 8'h00;
            15'd17102: data <= 8'h00;
            15'd17103: data <= 8'h00;
            15'd17104: data <= 8'h00;
            15'd17105: data <= 8'h03;
            15'd17106: data <= 8'hFF;
            15'd17107: data <= 8'hFF;
            15'd17108: data <= 8'hFF;
            15'd17109: data <= 8'hFF;
            15'd17110: data <= 8'hFF;
            15'd17111: data <= 8'hFF;
            15'd17112: data <= 8'hFF;
            15'd17113: data <= 8'hFF;
            15'd17114: data <= 8'hFF;
            15'd17115: data <= 8'hE0;
            15'd17116: data <= 8'hFF;
            15'd17117: data <= 8'hFF;
            15'd17118: data <= 8'hFF;
            15'd17119: data <= 8'hFF;
            15'd17120: data <= 8'hFF;
            15'd17121: data <= 8'hFF;
            15'd17122: data <= 8'hFF;
            15'd17123: data <= 8'hFF;
            15'd17124: data <= 8'h80;
            15'd17125: data <= 8'h00;
            15'd17126: data <= 8'h00;
            15'd17127: data <= 8'h00;
            15'd17128: data <= 8'h00;
            15'd17129: data <= 8'h00;
            15'd17130: data <= 8'h00;
            15'd17131: data <= 8'h00;
            15'd17132: data <= 8'h00;
            15'd17133: data <= 8'h00;
            15'd17134: data <= 8'h00;
            15'd17135: data <= 8'h03;
            15'd17136: data <= 8'hFF;
            15'd17137: data <= 8'hFF;
            15'd17138: data <= 8'hFF;
            15'd17139: data <= 8'hFF;
            15'd17140: data <= 8'hFF;
            15'd17141: data <= 8'hFF;
            15'd17142: data <= 8'hFF;
            15'd17143: data <= 8'hFF;
            15'd17144: data <= 8'hFF;
            15'd17145: data <= 8'h80;
            15'd17146: data <= 8'h3F;
            15'd17147: data <= 8'hFF;
            15'd17148: data <= 8'hFF;
            15'd17149: data <= 8'hFF;
            15'd17150: data <= 8'hFF;
            15'd17151: data <= 8'hFF;
            15'd17152: data <= 8'hFF;
            15'd17153: data <= 8'hFF;
            15'd17154: data <= 8'h80;
            15'd17155: data <= 8'h00;
            15'd17156: data <= 8'h00;
            15'd17157: data <= 8'h00;
            15'd17158: data <= 8'h00;
            15'd17159: data <= 8'h00;
            15'd17160: data <= 8'h00;
            15'd17161: data <= 8'h00;
            15'd17162: data <= 8'h00;
            15'd17163: data <= 8'h00;
            15'd17164: data <= 8'h00;
            15'd17165: data <= 8'h03;
            15'd17166: data <= 8'hFF;
            15'd17167: data <= 8'hFF;
            15'd17168: data <= 8'hFF;
            15'd17169: data <= 8'hFF;
            15'd17170: data <= 8'hFF;
            15'd17171: data <= 8'hFF;
            15'd17172: data <= 8'hFF;
            15'd17173: data <= 8'hFF;
            15'd17174: data <= 8'h80;
            15'd17175: data <= 8'h00;
            15'd17176: data <= 8'h1F;
            15'd17177: data <= 8'hFF;
            15'd17178: data <= 8'hFF;
            15'd17179: data <= 8'hFF;
            15'd17180: data <= 8'hFF;
            15'd17181: data <= 8'hFF;
            15'd17182: data <= 8'hFF;
            15'd17183: data <= 8'hFF;
            15'd17184: data <= 8'h80;
            15'd17185: data <= 8'h00;
            15'd17186: data <= 8'h00;
            15'd17187: data <= 8'h00;
            15'd17188: data <= 8'h00;
            15'd17189: data <= 8'h00;
            15'd17190: data <= 8'h00;
            15'd17191: data <= 8'h00;
            15'd17192: data <= 8'h00;
            15'd17193: data <= 8'h00;
            15'd17194: data <= 8'h00;
            15'd17195: data <= 8'h03;
            15'd17196: data <= 8'hFF;
            15'd17197: data <= 8'hFF;
            15'd17198: data <= 8'hFF;
            15'd17199: data <= 8'hFF;
            15'd17200: data <= 8'hFF;
            15'd17201: data <= 8'hFF;
            15'd17202: data <= 8'hFF;
            15'd17203: data <= 8'h80;
            15'd17204: data <= 8'h00;
            15'd17205: data <= 8'h00;
            15'd17206: data <= 8'h1F;
            15'd17207: data <= 8'hFF;
            15'd17208: data <= 8'hFF;
            15'd17209: data <= 8'hFF;
            15'd17210: data <= 8'hFF;
            15'd17211: data <= 8'hFF;
            15'd17212: data <= 8'hFF;
            15'd17213: data <= 8'hFF;
            15'd17214: data <= 8'h80;
            15'd17215: data <= 8'h00;
            15'd17216: data <= 8'h00;
            15'd17217: data <= 8'h00;
            15'd17218: data <= 8'h00;
            15'd17219: data <= 8'h00;
            15'd17220: data <= 8'h00;
            15'd17221: data <= 8'h00;
            15'd17222: data <= 8'h00;
            15'd17223: data <= 8'h00;
            15'd17224: data <= 8'h00;
            15'd17225: data <= 8'h03;
            15'd17226: data <= 8'hFF;
            15'd17227: data <= 8'hFF;
            15'd17228: data <= 8'hFF;
            15'd17229: data <= 8'hFF;
            15'd17230: data <= 8'hFF;
            15'd17231: data <= 8'hFF;
            15'd17232: data <= 8'hFE;
            15'd17233: data <= 8'h00;
            15'd17234: data <= 8'h00;
            15'd17235: data <= 8'h00;
            15'd17236: data <= 8'h1F;
            15'd17237: data <= 8'hFF;
            15'd17238: data <= 8'hFF;
            15'd17239: data <= 8'hFF;
            15'd17240: data <= 8'hFF;
            15'd17241: data <= 8'hFF;
            15'd17242: data <= 8'hFF;
            15'd17243: data <= 8'hFF;
            15'd17244: data <= 8'h80;
            15'd17245: data <= 8'h00;
            15'd17246: data <= 8'h00;
            15'd17247: data <= 8'h00;
            15'd17248: data <= 8'h00;
            15'd17249: data <= 8'h00;
            15'd17250: data <= 8'h00;
            15'd17251: data <= 8'h00;
            15'd17252: data <= 8'h00;
            15'd17253: data <= 8'h00;
            15'd17254: data <= 8'h00;
            15'd17255: data <= 8'h03;
            15'd17256: data <= 8'hFF;
            15'd17257: data <= 8'hFF;
            15'd17258: data <= 8'hFF;
            15'd17259: data <= 8'hFF;
            15'd17260: data <= 8'hFF;
            15'd17261: data <= 8'hFF;
            15'd17262: data <= 8'h80;
            15'd17263: data <= 8'h00;
            15'd17264: data <= 8'h00;
            15'd17265: data <= 8'h00;
            15'd17266: data <= 8'h0F;
            15'd17267: data <= 8'hFF;
            15'd17268: data <= 8'hFF;
            15'd17269: data <= 8'hFF;
            15'd17270: data <= 8'hFF;
            15'd17271: data <= 8'hFF;
            15'd17272: data <= 8'hFF;
            15'd17273: data <= 8'hFF;
            15'd17274: data <= 8'h80;
            15'd17275: data <= 8'h00;
            15'd17276: data <= 8'h00;
            15'd17277: data <= 8'h00;
            15'd17278: data <= 8'h00;
            15'd17279: data <= 8'h00;
            15'd17280: data <= 8'h00;
            15'd17281: data <= 8'h00;
            15'd17282: data <= 8'h00;
            15'd17283: data <= 8'h00;
            15'd17284: data <= 8'h00;
            15'd17285: data <= 8'h03;
            15'd17286: data <= 8'hFF;
            15'd17287: data <= 8'hFF;
            15'd17288: data <= 8'hFF;
            15'd17289: data <= 8'hFF;
            15'd17290: data <= 8'hFF;
            15'd17291: data <= 8'hFE;
            15'd17292: data <= 8'h00;
            15'd17293: data <= 8'h00;
            15'd17294: data <= 8'h00;
            15'd17295: data <= 8'h00;
            15'd17296: data <= 8'h07;
            15'd17297: data <= 8'hFF;
            15'd17298: data <= 8'hFF;
            15'd17299: data <= 8'hFF;
            15'd17300: data <= 8'hFF;
            15'd17301: data <= 8'hFF;
            15'd17302: data <= 8'hFF;
            15'd17303: data <= 8'hFF;
            15'd17304: data <= 8'h80;
            15'd17305: data <= 8'h00;
            15'd17306: data <= 8'h00;
            15'd17307: data <= 8'h00;
            15'd17308: data <= 8'h00;
            15'd17309: data <= 8'h00;
            15'd17310: data <= 8'h00;
            15'd17311: data <= 8'h00;
            15'd17312: data <= 8'h00;
            15'd17313: data <= 8'h00;
            15'd17314: data <= 8'h00;
            15'd17315: data <= 8'h03;
            15'd17316: data <= 8'hFF;
            15'd17317: data <= 8'hFF;
            15'd17318: data <= 8'hFF;
            15'd17319: data <= 8'hFF;
            15'd17320: data <= 8'hFF;
            15'd17321: data <= 8'hF0;
            15'd17322: data <= 8'h00;
            15'd17323: data <= 8'h00;
            15'd17324: data <= 8'h00;
            15'd17325: data <= 8'h10;
            15'd17326: data <= 8'h07;
            15'd17327: data <= 8'hFF;
            15'd17328: data <= 8'hFF;
            15'd17329: data <= 8'hFF;
            15'd17330: data <= 8'hFF;
            15'd17331: data <= 8'hFF;
            15'd17332: data <= 8'hFF;
            15'd17333: data <= 8'hFF;
            15'd17334: data <= 8'h80;
            15'd17335: data <= 8'h00;
            15'd17336: data <= 8'h00;
            15'd17337: data <= 8'h00;
            15'd17338: data <= 8'h00;
            15'd17339: data <= 8'h00;
            15'd17340: data <= 8'h00;
            15'd17341: data <= 8'h00;
            15'd17342: data <= 8'h00;
            15'd17343: data <= 8'h00;
            15'd17344: data <= 8'h00;
            15'd17345: data <= 8'h03;
            15'd17346: data <= 8'hFF;
            15'd17347: data <= 8'hFF;
            15'd17348: data <= 8'hFF;
            15'd17349: data <= 8'hFF;
            15'd17350: data <= 8'hFF;
            15'd17351: data <= 8'hC0;
            15'd17352: data <= 8'h00;
            15'd17353: data <= 8'h00;
            15'd17354: data <= 8'h01;
            15'd17355: data <= 8'hFC;
            15'd17356: data <= 8'h03;
            15'd17357: data <= 8'hFF;
            15'd17358: data <= 8'hFF;
            15'd17359: data <= 8'hFF;
            15'd17360: data <= 8'hFF;
            15'd17361: data <= 8'hFF;
            15'd17362: data <= 8'hFF;
            15'd17363: data <= 8'hFF;
            15'd17364: data <= 8'h80;
            15'd17365: data <= 8'h00;
            15'd17366: data <= 8'h00;
            15'd17367: data <= 8'h00;
            15'd17368: data <= 8'h00;
            15'd17369: data <= 8'h00;
            15'd17370: data <= 8'h00;
            15'd17371: data <= 8'h00;
            15'd17372: data <= 8'h00;
            15'd17373: data <= 8'h00;
            15'd17374: data <= 8'h00;
            15'd17375: data <= 8'h03;
            15'd17376: data <= 8'hFF;
            15'd17377: data <= 8'hFF;
            15'd17378: data <= 8'hFF;
            15'd17379: data <= 8'hFF;
            15'd17380: data <= 8'hFE;
            15'd17381: data <= 8'h00;
            15'd17382: data <= 8'h00;
            15'd17383: data <= 8'h00;
            15'd17384: data <= 8'hFF;
            15'd17385: data <= 8'hFE;
            15'd17386: data <= 8'h00;
            15'd17387: data <= 8'h7F;
            15'd17388: data <= 8'hFF;
            15'd17389: data <= 8'hFF;
            15'd17390: data <= 8'hFF;
            15'd17391: data <= 8'hFF;
            15'd17392: data <= 8'hFF;
            15'd17393: data <= 8'hFF;
            15'd17394: data <= 8'h80;
            15'd17395: data <= 8'h00;
            15'd17396: data <= 8'h00;
            15'd17397: data <= 8'h00;
            15'd17398: data <= 8'h00;
            15'd17399: data <= 8'h00;
            15'd17400: data <= 8'h00;
            15'd17401: data <= 8'h00;
            15'd17402: data <= 8'h00;
            15'd17403: data <= 8'h00;
            15'd17404: data <= 8'h00;
            15'd17405: data <= 8'h03;
            15'd17406: data <= 8'hFF;
            15'd17407: data <= 8'hFF;
            15'd17408: data <= 8'hFF;
            15'd17409: data <= 8'hFF;
            15'd17410: data <= 8'hF8;
            15'd17411: data <= 8'h00;
            15'd17412: data <= 8'h00;
            15'd17413: data <= 8'h3F;
            15'd17414: data <= 8'hFF;
            15'd17415: data <= 8'hFE;
            15'd17416: data <= 8'h00;
            15'd17417: data <= 8'h1F;
            15'd17418: data <= 8'hFF;
            15'd17419: data <= 8'hFF;
            15'd17420: data <= 8'hFF;
            15'd17421: data <= 8'hFF;
            15'd17422: data <= 8'hFF;
            15'd17423: data <= 8'hFF;
            15'd17424: data <= 8'h80;
            15'd17425: data <= 8'h00;
            15'd17426: data <= 8'h00;
            15'd17427: data <= 8'h00;
            15'd17428: data <= 8'h00;
            15'd17429: data <= 8'h00;
            15'd17430: data <= 8'h00;
            15'd17431: data <= 8'h00;
            15'd17432: data <= 8'h00;
            15'd17433: data <= 8'h00;
            15'd17434: data <= 8'h00;
            15'd17435: data <= 8'h03;
            15'd17436: data <= 8'hFF;
            15'd17437: data <= 8'hFF;
            15'd17438: data <= 8'hFF;
            15'd17439: data <= 8'hFF;
            15'd17440: data <= 8'hC0;
            15'd17441: data <= 8'h00;
            15'd17442: data <= 8'h07;
            15'd17443: data <= 8'hFF;
            15'd17444: data <= 8'hFF;
            15'd17445: data <= 8'hFF;
            15'd17446: data <= 8'h00;
            15'd17447: data <= 8'h03;
            15'd17448: data <= 8'hFF;
            15'd17449: data <= 8'hFF;
            15'd17450: data <= 8'hFF;
            15'd17451: data <= 8'hFF;
            15'd17452: data <= 8'hFF;
            15'd17453: data <= 8'hFF;
            15'd17454: data <= 8'h80;
            15'd17455: data <= 8'h00;
            15'd17456: data <= 8'h00;
            15'd17457: data <= 8'h00;
            15'd17458: data <= 8'h00;
            15'd17459: data <= 8'h00;
            15'd17460: data <= 8'h00;
            15'd17461: data <= 8'h00;
            15'd17462: data <= 8'h00;
            15'd17463: data <= 8'h00;
            15'd17464: data <= 8'h00;
            15'd17465: data <= 8'h03;
            15'd17466: data <= 8'hFF;
            15'd17467: data <= 8'hFF;
            15'd17468: data <= 8'hFF;
            15'd17469: data <= 8'hFF;
            15'd17470: data <= 8'h00;
            15'd17471: data <= 8'h00;
            15'd17472: data <= 8'h3F;
            15'd17473: data <= 8'hFF;
            15'd17474: data <= 8'hFF;
            15'd17475: data <= 8'hFF;
            15'd17476: data <= 8'h80;
            15'd17477: data <= 8'h00;
            15'd17478: data <= 8'h7F;
            15'd17479: data <= 8'hFF;
            15'd17480: data <= 8'hFF;
            15'd17481: data <= 8'hFF;
            15'd17482: data <= 8'hFF;
            15'd17483: data <= 8'hFF;
            15'd17484: data <= 8'h80;
            15'd17485: data <= 8'h00;
            15'd17486: data <= 8'h00;
            15'd17487: data <= 8'h00;
            15'd17488: data <= 8'h00;
            15'd17489: data <= 8'h00;
            15'd17490: data <= 8'h00;
            15'd17491: data <= 8'h00;
            15'd17492: data <= 8'h00;
            15'd17493: data <= 8'h00;
            15'd17494: data <= 8'h00;
            15'd17495: data <= 8'h03;
            15'd17496: data <= 8'hFF;
            15'd17497: data <= 8'hFF;
            15'd17498: data <= 8'hFF;
            15'd17499: data <= 8'hFE;
            15'd17500: data <= 8'h00;
            15'd17501: data <= 8'h01;
            15'd17502: data <= 8'hFF;
            15'd17503: data <= 8'hFF;
            15'd17504: data <= 8'hFF;
            15'd17505: data <= 8'hFF;
            15'd17506: data <= 8'hC0;
            15'd17507: data <= 8'h00;
            15'd17508: data <= 8'h04;
            15'd17509: data <= 8'h03;
            15'd17510: data <= 8'hFF;
            15'd17511: data <= 8'hFF;
            15'd17512: data <= 8'hFF;
            15'd17513: data <= 8'hFF;
            15'd17514: data <= 8'h80;
            15'd17515: data <= 8'h00;
            15'd17516: data <= 8'h00;
            15'd17517: data <= 8'h00;
            15'd17518: data <= 8'h00;
            15'd17519: data <= 8'h00;
            15'd17520: data <= 8'h00;
            15'd17521: data <= 8'h00;
            15'd17522: data <= 8'h00;
            15'd17523: data <= 8'h00;
            15'd17524: data <= 8'h00;
            15'd17525: data <= 8'h03;
            15'd17526: data <= 8'hFF;
            15'd17527: data <= 8'hFF;
            15'd17528: data <= 8'hFF;
            15'd17529: data <= 8'hFC;
            15'd17530: data <= 8'h00;
            15'd17531: data <= 8'h0F;
            15'd17532: data <= 8'hFF;
            15'd17533: data <= 8'hFF;
            15'd17534: data <= 8'hFF;
            15'd17535: data <= 8'hFF;
            15'd17536: data <= 8'hF0;
            15'd17537: data <= 8'h00;
            15'd17538: data <= 8'h00;
            15'd17539: data <= 8'h01;
            15'd17540: data <= 8'hFF;
            15'd17541: data <= 8'hFF;
            15'd17542: data <= 8'hFF;
            15'd17543: data <= 8'hFF;
            15'd17544: data <= 8'h80;
            15'd17545: data <= 8'h00;
            15'd17546: data <= 8'h00;
            15'd17547: data <= 8'h00;
            15'd17548: data <= 8'h00;
            15'd17549: data <= 8'h00;
            15'd17550: data <= 8'h00;
            15'd17551: data <= 8'h00;
            15'd17552: data <= 8'h00;
            15'd17553: data <= 8'h00;
            15'd17554: data <= 8'h00;
            15'd17555: data <= 8'h03;
            15'd17556: data <= 8'hFF;
            15'd17557: data <= 8'hFF;
            15'd17558: data <= 8'hFF;
            15'd17559: data <= 8'hF0;
            15'd17560: data <= 8'h00;
            15'd17561: data <= 8'h7F;
            15'd17562: data <= 8'hFF;
            15'd17563: data <= 8'hFF;
            15'd17564: data <= 8'hFF;
            15'd17565: data <= 8'hFF;
            15'd17566: data <= 8'hFC;
            15'd17567: data <= 8'h00;
            15'd17568: data <= 8'h00;
            15'd17569: data <= 8'h00;
            15'd17570: data <= 8'hFF;
            15'd17571: data <= 8'hFF;
            15'd17572: data <= 8'hFF;
            15'd17573: data <= 8'hFF;
            15'd17574: data <= 8'h80;
            15'd17575: data <= 8'h00;
            15'd17576: data <= 8'h00;
            15'd17577: data <= 8'h00;
            15'd17578: data <= 8'h00;
            15'd17579: data <= 8'h00;
            15'd17580: data <= 8'h00;
            15'd17581: data <= 8'h00;
            15'd17582: data <= 8'h00;
            15'd17583: data <= 8'h00;
            15'd17584: data <= 8'h00;
            15'd17585: data <= 8'h03;
            15'd17586: data <= 8'hFF;
            15'd17587: data <= 8'hFF;
            15'd17588: data <= 8'hFF;
            15'd17589: data <= 8'hE0;
            15'd17590: data <= 8'h03;
            15'd17591: data <= 8'hFF;
            15'd17592: data <= 8'hFF;
            15'd17593: data <= 8'hFF;
            15'd17594: data <= 8'hFF;
            15'd17595: data <= 8'hFF;
            15'd17596: data <= 8'hFF;
            15'd17597: data <= 8'h00;
            15'd17598: data <= 8'h00;
            15'd17599: data <= 8'h00;
            15'd17600: data <= 8'h7F;
            15'd17601: data <= 8'hFF;
            15'd17602: data <= 8'hFF;
            15'd17603: data <= 8'hFF;
            15'd17604: data <= 8'h80;
            15'd17605: data <= 8'h00;
            15'd17606: data <= 8'h00;
            15'd17607: data <= 8'h00;
            15'd17608: data <= 8'h00;
            15'd17609: data <= 8'h00;
            15'd17610: data <= 8'h00;
            15'd17611: data <= 8'h00;
            15'd17612: data <= 8'h00;
            15'd17613: data <= 8'h00;
            15'd17614: data <= 8'h00;
            15'd17615: data <= 8'h03;
            15'd17616: data <= 8'hFF;
            15'd17617: data <= 8'hFF;
            15'd17618: data <= 8'hFF;
            15'd17619: data <= 8'h80;
            15'd17620: data <= 8'h07;
            15'd17621: data <= 8'hFF;
            15'd17622: data <= 8'hFF;
            15'd17623: data <= 8'hFF;
            15'd17624: data <= 8'hFF;
            15'd17625: data <= 8'hFF;
            15'd17626: data <= 8'hFF;
            15'd17627: data <= 8'hE0;
            15'd17628: data <= 8'h00;
            15'd17629: data <= 8'h00;
            15'd17630: data <= 8'h7F;
            15'd17631: data <= 8'hFF;
            15'd17632: data <= 8'hFF;
            15'd17633: data <= 8'hFF;
            15'd17634: data <= 8'h80;
            15'd17635: data <= 8'h00;
            15'd17636: data <= 8'h00;
            15'd17637: data <= 8'h00;
            15'd17638: data <= 8'h00;
            15'd17639: data <= 8'h00;
            15'd17640: data <= 8'h00;
            15'd17641: data <= 8'h00;
            15'd17642: data <= 8'h00;
            15'd17643: data <= 8'h00;
            15'd17644: data <= 8'h00;
            15'd17645: data <= 8'h03;
            15'd17646: data <= 8'hFF;
            15'd17647: data <= 8'hFF;
            15'd17648: data <= 8'hFF;
            15'd17649: data <= 8'h00;
            15'd17650: data <= 8'h0F;
            15'd17651: data <= 8'hFF;
            15'd17652: data <= 8'hFF;
            15'd17653: data <= 8'hFF;
            15'd17654: data <= 8'hFF;
            15'd17655: data <= 8'hFF;
            15'd17656: data <= 8'hFF;
            15'd17657: data <= 8'hFE;
            15'd17658: data <= 8'h00;
            15'd17659: data <= 8'h00;
            15'd17660: data <= 8'h3F;
            15'd17661: data <= 8'hFF;
            15'd17662: data <= 8'hFF;
            15'd17663: data <= 8'hFF;
            15'd17664: data <= 8'h80;
            15'd17665: data <= 8'h00;
            15'd17666: data <= 8'h00;
            15'd17667: data <= 8'h00;
            15'd17668: data <= 8'h00;
            15'd17669: data <= 8'h00;
            15'd17670: data <= 8'h00;
            15'd17671: data <= 8'h00;
            15'd17672: data <= 8'h00;
            15'd17673: data <= 8'h00;
            15'd17674: data <= 8'h00;
            15'd17675: data <= 8'h03;
            15'd17676: data <= 8'hFF;
            15'd17677: data <= 8'hFF;
            15'd17678: data <= 8'hFE;
            15'd17679: data <= 8'h00;
            15'd17680: data <= 8'h3F;
            15'd17681: data <= 8'hFF;
            15'd17682: data <= 8'hFF;
            15'd17683: data <= 8'hFF;
            15'd17684: data <= 8'hFF;
            15'd17685: data <= 8'hFF;
            15'd17686: data <= 8'hFF;
            15'd17687: data <= 8'hFF;
            15'd17688: data <= 8'h80;
            15'd17689: data <= 8'h00;
            15'd17690: data <= 8'h3F;
            15'd17691: data <= 8'hFF;
            15'd17692: data <= 8'hFF;
            15'd17693: data <= 8'hFF;
            15'd17694: data <= 8'h80;
            15'd17695: data <= 8'h00;
            15'd17696: data <= 8'h00;
            15'd17697: data <= 8'h00;
            15'd17698: data <= 8'h00;
            15'd17699: data <= 8'h00;
            15'd17700: data <= 8'h00;
            15'd17701: data <= 8'h00;
            15'd17702: data <= 8'h00;
            15'd17703: data <= 8'h00;
            15'd17704: data <= 8'h00;
            15'd17705: data <= 8'h03;
            15'd17706: data <= 8'hFF;
            15'd17707: data <= 8'hFF;
            15'd17708: data <= 8'hFC;
            15'd17709: data <= 8'h00;
            15'd17710: data <= 8'hFF;
            15'd17711: data <= 8'hFF;
            15'd17712: data <= 8'hFF;
            15'd17713: data <= 8'hFF;
            15'd17714: data <= 8'hFF;
            15'd17715: data <= 8'hFF;
            15'd17716: data <= 8'hFF;
            15'd17717: data <= 8'hFF;
            15'd17718: data <= 8'hFF;
            15'd17719: data <= 8'hE0;
            15'd17720: data <= 8'h3F;
            15'd17721: data <= 8'hFF;
            15'd17722: data <= 8'hFF;
            15'd17723: data <= 8'hFF;
            15'd17724: data <= 8'h80;
            15'd17725: data <= 8'h00;
            15'd17726: data <= 8'h00;
            15'd17727: data <= 8'h00;
            15'd17728: data <= 8'h00;
            15'd17729: data <= 8'h00;
            15'd17730: data <= 8'h00;
            15'd17731: data <= 8'h00;
            15'd17732: data <= 8'h00;
            15'd17733: data <= 8'h00;
            15'd17734: data <= 8'h00;
            15'd17735: data <= 8'h03;
            15'd17736: data <= 8'hFF;
            15'd17737: data <= 8'hFF;
            15'd17738: data <= 8'hF8;
            15'd17739: data <= 8'h01;
            15'd17740: data <= 8'hFF;
            15'd17741: data <= 8'hFF;
            15'd17742: data <= 8'hFF;
            15'd17743: data <= 8'hFF;
            15'd17744: data <= 8'hFF;
            15'd17745: data <= 8'hFF;
            15'd17746: data <= 8'hFF;
            15'd17747: data <= 8'hFF;
            15'd17748: data <= 8'hFF;
            15'd17749: data <= 8'hF0;
            15'd17750: data <= 8'h1F;
            15'd17751: data <= 8'hFF;
            15'd17752: data <= 8'hFF;
            15'd17753: data <= 8'hFF;
            15'd17754: data <= 8'h80;
            15'd17755: data <= 8'h00;
            15'd17756: data <= 8'h00;
            15'd17757: data <= 8'h00;
            15'd17758: data <= 8'h00;
            15'd17759: data <= 8'h00;
            15'd17760: data <= 8'h00;
            15'd17761: data <= 8'h00;
            15'd17762: data <= 8'h00;
            15'd17763: data <= 8'h00;
            15'd17764: data <= 8'h00;
            15'd17765: data <= 8'h03;
            15'd17766: data <= 8'hFF;
            15'd17767: data <= 8'hFF;
            15'd17768: data <= 8'hF0;
            15'd17769: data <= 8'h03;
            15'd17770: data <= 8'hFF;
            15'd17771: data <= 8'hFF;
            15'd17772: data <= 8'hFF;
            15'd17773: data <= 8'hFF;
            15'd17774: data <= 8'hFF;
            15'd17775: data <= 8'hFF;
            15'd17776: data <= 8'hFF;
            15'd17777: data <= 8'hFF;
            15'd17778: data <= 8'hFF;
            15'd17779: data <= 8'hF0;
            15'd17780: data <= 8'h1F;
            15'd17781: data <= 8'hFF;
            15'd17782: data <= 8'hFF;
            15'd17783: data <= 8'hFF;
            15'd17784: data <= 8'h80;
            15'd17785: data <= 8'h00;
            15'd17786: data <= 8'h00;
            15'd17787: data <= 8'h00;
            15'd17788: data <= 8'h00;
            15'd17789: data <= 8'h00;
            15'd17790: data <= 8'h00;
            15'd17791: data <= 8'h00;
            15'd17792: data <= 8'h00;
            15'd17793: data <= 8'h00;
            15'd17794: data <= 8'h00;
            15'd17795: data <= 8'h03;
            15'd17796: data <= 8'hFF;
            15'd17797: data <= 8'hFF;
            15'd17798: data <= 8'hF0;
            15'd17799: data <= 8'h0F;
            15'd17800: data <= 8'hFF;
            15'd17801: data <= 8'hFF;
            15'd17802: data <= 8'hFF;
            15'd17803: data <= 8'hFF;
            15'd17804: data <= 8'hFF;
            15'd17805: data <= 8'hFF;
            15'd17806: data <= 8'hFF;
            15'd17807: data <= 8'hFF;
            15'd17808: data <= 8'hFF;
            15'd17809: data <= 8'hF0;
            15'd17810: data <= 8'h1F;
            15'd17811: data <= 8'hFF;
            15'd17812: data <= 8'hFF;
            15'd17813: data <= 8'hFF;
            15'd17814: data <= 8'h80;
            15'd17815: data <= 8'h00;
            15'd17816: data <= 8'h00;
            15'd17817: data <= 8'h00;
            15'd17818: data <= 8'h00;
            15'd17819: data <= 8'h00;
            15'd17820: data <= 8'h00;
            15'd17821: data <= 8'h00;
            15'd17822: data <= 8'h00;
            15'd17823: data <= 8'h00;
            15'd17824: data <= 8'h00;
            15'd17825: data <= 8'h03;
            15'd17826: data <= 8'hFF;
            15'd17827: data <= 8'hFF;
            15'd17828: data <= 8'hE0;
            15'd17829: data <= 8'h0F;
            15'd17830: data <= 8'hFF;
            15'd17831: data <= 8'hFF;
            15'd17832: data <= 8'hFF;
            15'd17833: data <= 8'hFF;
            15'd17834: data <= 8'hFF;
            15'd17835: data <= 8'hFF;
            15'd17836: data <= 8'hFF;
            15'd17837: data <= 8'hFF;
            15'd17838: data <= 8'hFF;
            15'd17839: data <= 8'hF8;
            15'd17840: data <= 8'h0F;
            15'd17841: data <= 8'hFF;
            15'd17842: data <= 8'hFF;
            15'd17843: data <= 8'hFF;
            15'd17844: data <= 8'h80;
            15'd17845: data <= 8'h00;
            15'd17846: data <= 8'h00;
            15'd17847: data <= 8'h00;
            15'd17848: data <= 8'h00;
            15'd17849: data <= 8'h00;
            15'd17850: data <= 8'h00;
            15'd17851: data <= 8'h00;
            15'd17852: data <= 8'h00;
            15'd17853: data <= 8'h00;
            15'd17854: data <= 8'h00;
            15'd17855: data <= 8'h03;
            15'd17856: data <= 8'hFF;
            15'd17857: data <= 8'hFF;
            15'd17858: data <= 8'hC0;
            15'd17859: data <= 8'h1F;
            15'd17860: data <= 8'hFF;
            15'd17861: data <= 8'hFF;
            15'd17862: data <= 8'hFF;
            15'd17863: data <= 8'hFF;
            15'd17864: data <= 8'hFF;
            15'd17865: data <= 8'hFF;
            15'd17866: data <= 8'hFF;
            15'd17867: data <= 8'hFF;
            15'd17868: data <= 8'hFF;
            15'd17869: data <= 8'hF8;
            15'd17870: data <= 8'h0F;
            15'd17871: data <= 8'hFF;
            15'd17872: data <= 8'hFF;
            15'd17873: data <= 8'hFF;
            15'd17874: data <= 8'h80;
            15'd17875: data <= 8'h00;
            15'd17876: data <= 8'h00;
            15'd17877: data <= 8'h00;
            15'd17878: data <= 8'h00;
            15'd17879: data <= 8'h00;
            15'd17880: data <= 8'h00;
            15'd17881: data <= 8'h00;
            15'd17882: data <= 8'h00;
            15'd17883: data <= 8'h00;
            15'd17884: data <= 8'h00;
            15'd17885: data <= 8'h03;
            15'd17886: data <= 8'hFF;
            15'd17887: data <= 8'hFF;
            15'd17888: data <= 8'hC0;
            15'd17889: data <= 8'h7F;
            15'd17890: data <= 8'hFF;
            15'd17891: data <= 8'hFF;
            15'd17892: data <= 8'hFF;
            15'd17893: data <= 8'hFF;
            15'd17894: data <= 8'hFF;
            15'd17895: data <= 8'hFF;
            15'd17896: data <= 8'hFF;
            15'd17897: data <= 8'hFF;
            15'd17898: data <= 8'hFF;
            15'd17899: data <= 8'hF8;
            15'd17900: data <= 8'h0F;
            15'd17901: data <= 8'hFF;
            15'd17902: data <= 8'hFF;
            15'd17903: data <= 8'hFF;
            15'd17904: data <= 8'h80;
            15'd17905: data <= 8'h00;
            15'd17906: data <= 8'h00;
            15'd17907: data <= 8'h00;
            15'd17908: data <= 8'h00;
            15'd17909: data <= 8'h00;
            15'd17910: data <= 8'h00;
            15'd17911: data <= 8'h00;
            15'd17912: data <= 8'h00;
            15'd17913: data <= 8'h00;
            15'd17914: data <= 8'h00;
            15'd17915: data <= 8'h03;
            15'd17916: data <= 8'hFF;
            15'd17917: data <= 8'hFF;
            15'd17918: data <= 8'h80;
            15'd17919: data <= 8'h7F;
            15'd17920: data <= 8'hFF;
            15'd17921: data <= 8'hFF;
            15'd17922: data <= 8'hFF;
            15'd17923: data <= 8'hFF;
            15'd17924: data <= 8'hFF;
            15'd17925: data <= 8'hFF;
            15'd17926: data <= 8'hFF;
            15'd17927: data <= 8'hFF;
            15'd17928: data <= 8'hFF;
            15'd17929: data <= 8'hF8;
            15'd17930: data <= 8'h07;
            15'd17931: data <= 8'hFF;
            15'd17932: data <= 8'hFF;
            15'd17933: data <= 8'hFF;
            15'd17934: data <= 8'h80;
            15'd17935: data <= 8'h00;
            15'd17936: data <= 8'h00;
            15'd17937: data <= 8'h00;
            15'd17938: data <= 8'h00;
            15'd17939: data <= 8'h00;
            15'd17940: data <= 8'h00;
            15'd17941: data <= 8'h00;
            15'd17942: data <= 8'h00;
            15'd17943: data <= 8'h00;
            15'd17944: data <= 8'h00;
            15'd17945: data <= 8'h03;
            15'd17946: data <= 8'hFF;
            15'd17947: data <= 8'hFF;
            15'd17948: data <= 8'h80;
            15'd17949: data <= 8'hFF;
            15'd17950: data <= 8'hFF;
            15'd17951: data <= 8'hFF;
            15'd17952: data <= 8'hFF;
            15'd17953: data <= 8'hFF;
            15'd17954: data <= 8'hFF;
            15'd17955: data <= 8'hFF;
            15'd17956: data <= 8'hFF;
            15'd17957: data <= 8'hFF;
            15'd17958: data <= 8'hFF;
            15'd17959: data <= 8'hFC;
            15'd17960: data <= 8'h07;
            15'd17961: data <= 8'hFF;
            15'd17962: data <= 8'hFF;
            15'd17963: data <= 8'hFF;
            15'd17964: data <= 8'h80;
            15'd17965: data <= 8'h00;
            15'd17966: data <= 8'h00;
            15'd17967: data <= 8'h00;
            15'd17968: data <= 8'h00;
            15'd17969: data <= 8'h00;
            15'd17970: data <= 8'h00;
            15'd17971: data <= 8'h00;
            15'd17972: data <= 8'h00;
            15'd17973: data <= 8'h00;
            15'd17974: data <= 8'h00;
            15'd17975: data <= 8'h03;
            15'd17976: data <= 8'hFF;
            15'd17977: data <= 8'hFF;
            15'd17978: data <= 8'h00;
            15'd17979: data <= 8'hFF;
            15'd17980: data <= 8'hFF;
            15'd17981: data <= 8'hFF;
            15'd17982: data <= 8'hFF;
            15'd17983: data <= 8'hFF;
            15'd17984: data <= 8'hFF;
            15'd17985: data <= 8'hFF;
            15'd17986: data <= 8'hFF;
            15'd17987: data <= 8'hFF;
            15'd17988: data <= 8'hFF;
            15'd17989: data <= 8'hFC;
            15'd17990: data <= 8'h07;
            15'd17991: data <= 8'hFF;
            15'd17992: data <= 8'hFF;
            15'd17993: data <= 8'hFF;
            15'd17994: data <= 8'h80;
            15'd17995: data <= 8'h00;
            15'd17996: data <= 8'h00;
            15'd17997: data <= 8'h00;
            15'd17998: data <= 8'h00;
            15'd17999: data <= 8'h00;
            15'd18000: data <= 8'h00;
            15'd18001: data <= 8'h00;
            15'd18002: data <= 8'h00;
            15'd18003: data <= 8'h00;
            15'd18004: data <= 8'h00;
            15'd18005: data <= 8'h03;
            15'd18006: data <= 8'hFF;
            15'd18007: data <= 8'hFF;
            15'd18008: data <= 8'h01;
            15'd18009: data <= 8'hFF;
            15'd18010: data <= 8'hFF;
            15'd18011: data <= 8'hFF;
            15'd18012: data <= 8'hFF;
            15'd18013: data <= 8'hFF;
            15'd18014: data <= 8'hFF;
            15'd18015: data <= 8'hFF;
            15'd18016: data <= 8'hFF;
            15'd18017: data <= 8'hFF;
            15'd18018: data <= 8'hFF;
            15'd18019: data <= 8'hFE;
            15'd18020: data <= 8'h03;
            15'd18021: data <= 8'hFF;
            15'd18022: data <= 8'hFF;
            15'd18023: data <= 8'hFF;
            15'd18024: data <= 8'h80;
            15'd18025: data <= 8'h00;
            15'd18026: data <= 8'h00;
            15'd18027: data <= 8'h00;
            15'd18028: data <= 8'h00;
            15'd18029: data <= 8'h00;
            15'd18030: data <= 8'h00;
            15'd18031: data <= 8'h00;
            15'd18032: data <= 8'h00;
            15'd18033: data <= 8'h00;
            15'd18034: data <= 8'h00;
            15'd18035: data <= 8'h03;
            15'd18036: data <= 8'hFF;
            15'd18037: data <= 8'hFF;
            15'd18038: data <= 8'h01;
            15'd18039: data <= 8'hFF;
            15'd18040: data <= 8'hFF;
            15'd18041: data <= 8'hFF;
            15'd18042: data <= 8'hFF;
            15'd18043: data <= 8'hFF;
            15'd18044: data <= 8'hFF;
            15'd18045: data <= 8'hFF;
            15'd18046: data <= 8'hFF;
            15'd18047: data <= 8'hFF;
            15'd18048: data <= 8'hFF;
            15'd18049: data <= 8'hFE;
            15'd18050: data <= 8'h01;
            15'd18051: data <= 8'hFF;
            15'd18052: data <= 8'hFF;
            15'd18053: data <= 8'hFF;
            15'd18054: data <= 8'h80;
            15'd18055: data <= 8'h00;
            15'd18056: data <= 8'h00;
            15'd18057: data <= 8'h00;
            15'd18058: data <= 8'h00;
            15'd18059: data <= 8'h00;
            15'd18060: data <= 8'h00;
            15'd18061: data <= 8'h00;
            15'd18062: data <= 8'h00;
            15'd18063: data <= 8'h00;
            15'd18064: data <= 8'h00;
            15'd18065: data <= 8'h03;
            15'd18066: data <= 8'hFF;
            15'd18067: data <= 8'hFF;
            15'd18068: data <= 8'h01;
            15'd18069: data <= 8'hFF;
            15'd18070: data <= 8'hF9;
            15'd18071: data <= 8'hFF;
            15'd18072: data <= 8'hFF;
            15'd18073: data <= 8'hFF;
            15'd18074: data <= 8'hFF;
            15'd18075: data <= 8'hFF;
            15'd18076: data <= 8'hFF;
            15'd18077: data <= 8'hFF;
            15'd18078: data <= 8'hFF;
            15'd18079: data <= 8'hFE;
            15'd18080: data <= 8'h01;
            15'd18081: data <= 8'hFF;
            15'd18082: data <= 8'hFF;
            15'd18083: data <= 8'hFF;
            15'd18084: data <= 8'h80;
            15'd18085: data <= 8'h00;
            15'd18086: data <= 8'h00;
            15'd18087: data <= 8'h00;
            15'd18088: data <= 8'h00;
            15'd18089: data <= 8'h00;
            15'd18090: data <= 8'h00;
            15'd18091: data <= 8'h00;
            15'd18092: data <= 8'h00;
            15'd18093: data <= 8'h00;
            15'd18094: data <= 8'h00;
            15'd18095: data <= 8'h03;
            15'd18096: data <= 8'hFF;
            15'd18097: data <= 8'hFE;
            15'd18098: data <= 8'h03;
            15'd18099: data <= 8'hFF;
            15'd18100: data <= 8'hF0;
            15'd18101: data <= 8'hFF;
            15'd18102: data <= 8'hFF;
            15'd18103: data <= 8'hFF;
            15'd18104: data <= 8'hFF;
            15'd18105: data <= 8'hFF;
            15'd18106: data <= 8'hFF;
            15'd18107: data <= 8'hFF;
            15'd18108: data <= 8'hFF;
            15'd18109: data <= 8'hFF;
            15'd18110: data <= 8'h00;
            15'd18111: data <= 8'hFF;
            15'd18112: data <= 8'hFF;
            15'd18113: data <= 8'hFF;
            15'd18114: data <= 8'h80;
            15'd18115: data <= 8'h00;
            15'd18116: data <= 8'h00;
            15'd18117: data <= 8'h00;
            15'd18118: data <= 8'h00;
            15'd18119: data <= 8'h00;
            15'd18120: data <= 8'h00;
            15'd18121: data <= 8'h00;
            15'd18122: data <= 8'h00;
            15'd18123: data <= 8'h00;
            15'd18124: data <= 8'h00;
            15'd18125: data <= 8'h03;
            15'd18126: data <= 8'hFF;
            15'd18127: data <= 8'hFE;
            15'd18128: data <= 8'h03;
            15'd18129: data <= 8'hFF;
            15'd18130: data <= 8'hF0;
            15'd18131: data <= 8'hFF;
            15'd18132: data <= 8'hC7;
            15'd18133: data <= 8'hFF;
            15'd18134: data <= 8'hFF;
            15'd18135: data <= 8'hFF;
            15'd18136: data <= 8'hFF;
            15'd18137: data <= 8'hFF;
            15'd18138: data <= 8'hFF;
            15'd18139: data <= 8'hFF;
            15'd18140: data <= 8'h00;
            15'd18141: data <= 8'hFF;
            15'd18142: data <= 8'hFF;
            15'd18143: data <= 8'hFF;
            15'd18144: data <= 8'h80;
            15'd18145: data <= 8'h00;
            15'd18146: data <= 8'h00;
            15'd18147: data <= 8'h00;
            15'd18148: data <= 8'h00;
            15'd18149: data <= 8'h00;
            15'd18150: data <= 8'h00;
            15'd18151: data <= 8'h00;
            15'd18152: data <= 8'h00;
            15'd18153: data <= 8'h00;
            15'd18154: data <= 8'h00;
            15'd18155: data <= 8'h03;
            15'd18156: data <= 8'hFF;
            15'd18157: data <= 8'hFE;
            15'd18158: data <= 8'h07;
            15'd18159: data <= 8'hFF;
            15'd18160: data <= 8'hF0;
            15'd18161: data <= 8'hFF;
            15'd18162: data <= 8'h83;
            15'd18163: data <= 8'hFF;
            15'd18164: data <= 8'hFF;
            15'd18165: data <= 8'hFF;
            15'd18166: data <= 8'hFF;
            15'd18167: data <= 8'hFF;
            15'd18168: data <= 8'hFF;
            15'd18169: data <= 8'hFF;
            15'd18170: data <= 8'h80;
            15'd18171: data <= 8'h7F;
            15'd18172: data <= 8'hFF;
            15'd18173: data <= 8'hFF;
            15'd18174: data <= 8'h80;
            15'd18175: data <= 8'h00;
            15'd18176: data <= 8'h00;
            15'd18177: data <= 8'h00;
            15'd18178: data <= 8'h00;
            15'd18179: data <= 8'h00;
            15'd18180: data <= 8'h00;
            15'd18181: data <= 8'h00;
            15'd18182: data <= 8'h00;
            15'd18183: data <= 8'h00;
            15'd18184: data <= 8'h00;
            15'd18185: data <= 8'h03;
            15'd18186: data <= 8'hFF;
            15'd18187: data <= 8'hFE;
            15'd18188: data <= 8'h07;
            15'd18189: data <= 8'hFF;
            15'd18190: data <= 8'hFD;
            15'd18191: data <= 8'hFF;
            15'd18192: data <= 8'h83;
            15'd18193: data <= 8'hFF;
            15'd18194: data <= 8'hFF;
            15'd18195: data <= 8'hFF;
            15'd18196: data <= 8'hFF;
            15'd18197: data <= 8'hFF;
            15'd18198: data <= 8'hFF;
            15'd18199: data <= 8'hFF;
            15'd18200: data <= 8'h80;
            15'd18201: data <= 8'h7F;
            15'd18202: data <= 8'hFF;
            15'd18203: data <= 8'hFF;
            15'd18204: data <= 8'h80;
            15'd18205: data <= 8'h00;
            15'd18206: data <= 8'h00;
            15'd18207: data <= 8'h00;
            15'd18208: data <= 8'h00;
            15'd18209: data <= 8'h00;
            15'd18210: data <= 8'h00;
            15'd18211: data <= 8'h00;
            15'd18212: data <= 8'h00;
            15'd18213: data <= 8'h00;
            15'd18214: data <= 8'h00;
            15'd18215: data <= 8'h03;
            15'd18216: data <= 8'hFF;
            15'd18217: data <= 8'hFE;
            15'd18218: data <= 8'h07;
            15'd18219: data <= 8'hFF;
            15'd18220: data <= 8'hFF;
            15'd18221: data <= 8'hFF;
            15'd18222: data <= 8'h83;
            15'd18223: data <= 8'hFF;
            15'd18224: data <= 8'hFF;
            15'd18225: data <= 8'hFF;
            15'd18226: data <= 8'hFF;
            15'd18227: data <= 8'hFF;
            15'd18228: data <= 8'hFF;
            15'd18229: data <= 8'hFF;
            15'd18230: data <= 8'hC0;
            15'd18231: data <= 8'h3F;
            15'd18232: data <= 8'hFF;
            15'd18233: data <= 8'hFF;
            15'd18234: data <= 8'h80;
            15'd18235: data <= 8'h00;
            15'd18236: data <= 8'h00;
            15'd18237: data <= 8'h00;
            15'd18238: data <= 8'h00;
            15'd18239: data <= 8'h00;
            15'd18240: data <= 8'h00;
            15'd18241: data <= 8'h00;
            15'd18242: data <= 8'h00;
            15'd18243: data <= 8'h00;
            15'd18244: data <= 8'h00;
            15'd18245: data <= 8'h03;
            15'd18246: data <= 8'hFF;
            15'd18247: data <= 8'hFE;
            15'd18248: data <= 8'h07;
            15'd18249: data <= 8'hFF;
            15'd18250: data <= 8'hFF;
            15'd18251: data <= 8'hFF;
            15'd18252: data <= 8'hEF;
            15'd18253: data <= 8'hFF;
            15'd18254: data <= 8'hFF;
            15'd18255: data <= 8'hFF;
            15'd18256: data <= 8'hFF;
            15'd18257: data <= 8'hFF;
            15'd18258: data <= 8'hFF;
            15'd18259: data <= 8'hFF;
            15'd18260: data <= 8'hE0;
            15'd18261: data <= 8'h3F;
            15'd18262: data <= 8'hFF;
            15'd18263: data <= 8'hFF;
            15'd18264: data <= 8'h80;
            15'd18265: data <= 8'h00;
            15'd18266: data <= 8'h00;
            15'd18267: data <= 8'h00;
            15'd18268: data <= 8'h00;
            15'd18269: data <= 8'h00;
            15'd18270: data <= 8'h00;
            15'd18271: data <= 8'h00;
            15'd18272: data <= 8'h00;
            15'd18273: data <= 8'h00;
            15'd18274: data <= 8'h00;
            15'd18275: data <= 8'h03;
            15'd18276: data <= 8'hFF;
            15'd18277: data <= 8'hFE;
            15'd18278: data <= 8'h07;
            15'd18279: data <= 8'hFF;
            15'd18280: data <= 8'hFF;
            15'd18281: data <= 8'hFF;
            15'd18282: data <= 8'hFF;
            15'd18283: data <= 8'hFF;
            15'd18284: data <= 8'hFF;
            15'd18285: data <= 8'hFF;
            15'd18286: data <= 8'hFF;
            15'd18287: data <= 8'hFF;
            15'd18288: data <= 8'hFF;
            15'd18289: data <= 8'hFF;
            15'd18290: data <= 8'hE0;
            15'd18291: data <= 8'h1F;
            15'd18292: data <= 8'hFF;
            15'd18293: data <= 8'hFF;
            15'd18294: data <= 8'h80;
            15'd18295: data <= 8'h00;
            15'd18296: data <= 8'h00;
            15'd18297: data <= 8'h00;
            15'd18298: data <= 8'h00;
            15'd18299: data <= 8'h00;
            15'd18300: data <= 8'h00;
            15'd18301: data <= 8'h00;
            15'd18302: data <= 8'h00;
            15'd18303: data <= 8'h00;
            15'd18304: data <= 8'h00;
            15'd18305: data <= 8'h03;
            15'd18306: data <= 8'hFF;
            15'd18307: data <= 8'hFE;
            15'd18308: data <= 8'h07;
            15'd18309: data <= 8'hFF;
            15'd18310: data <= 8'hFF;
            15'd18311: data <= 8'hFF;
            15'd18312: data <= 8'hFF;
            15'd18313: data <= 8'hFF;
            15'd18314: data <= 8'hFF;
            15'd18315: data <= 8'hFF;
            15'd18316: data <= 8'hFF;
            15'd18317: data <= 8'hFF;
            15'd18318: data <= 8'hFF;
            15'd18319: data <= 8'hFF;
            15'd18320: data <= 8'hF0;
            15'd18321: data <= 8'h0F;
            15'd18322: data <= 8'hFF;
            15'd18323: data <= 8'hFF;
            15'd18324: data <= 8'h80;
            15'd18325: data <= 8'h00;
            15'd18326: data <= 8'h00;
            15'd18327: data <= 8'h00;
            15'd18328: data <= 8'h00;
            15'd18329: data <= 8'h00;
            15'd18330: data <= 8'h00;
            15'd18331: data <= 8'h00;
            15'd18332: data <= 8'h00;
            15'd18333: data <= 8'h00;
            15'd18334: data <= 8'h00;
            15'd18335: data <= 8'h03;
            15'd18336: data <= 8'hFF;
            15'd18337: data <= 8'hFE;
            15'd18338: data <= 8'h07;
            15'd18339: data <= 8'hFF;
            15'd18340: data <= 8'hFF;
            15'd18341: data <= 8'hFF;
            15'd18342: data <= 8'hFF;
            15'd18343: data <= 8'hFF;
            15'd18344: data <= 8'hFF;
            15'd18345: data <= 8'hFF;
            15'd18346: data <= 8'hFF;
            15'd18347: data <= 8'hFF;
            15'd18348: data <= 8'hFF;
            15'd18349: data <= 8'hFF;
            15'd18350: data <= 8'hF0;
            15'd18351: data <= 8'h0F;
            15'd18352: data <= 8'hFF;
            15'd18353: data <= 8'hFF;
            15'd18354: data <= 8'h80;
            15'd18355: data <= 8'h00;
            15'd18356: data <= 8'h00;
            15'd18357: data <= 8'h00;
            15'd18358: data <= 8'h00;
            15'd18359: data <= 8'h00;
            15'd18360: data <= 8'h00;
            15'd18361: data <= 8'h00;
            15'd18362: data <= 8'h00;
            15'd18363: data <= 8'h00;
            15'd18364: data <= 8'h00;
            15'd18365: data <= 8'h03;
            15'd18366: data <= 8'hFF;
            15'd18367: data <= 8'hFE;
            15'd18368: data <= 8'h07;
            15'd18369: data <= 8'hFF;
            15'd18370: data <= 8'hFF;
            15'd18371: data <= 8'hFF;
            15'd18372: data <= 8'hFF;
            15'd18373: data <= 8'hFF;
            15'd18374: data <= 8'hFF;
            15'd18375: data <= 8'hFF;
            15'd18376: data <= 8'hFF;
            15'd18377: data <= 8'hFF;
            15'd18378: data <= 8'hFF;
            15'd18379: data <= 8'hFF;
            15'd18380: data <= 8'hF8;
            15'd18381: data <= 8'h0F;
            15'd18382: data <= 8'hFF;
            15'd18383: data <= 8'hFF;
            15'd18384: data <= 8'h80;
            15'd18385: data <= 8'h00;
            15'd18386: data <= 8'h00;
            15'd18387: data <= 8'h00;
            15'd18388: data <= 8'h00;
            15'd18389: data <= 8'h00;
            15'd18390: data <= 8'h00;
            15'd18391: data <= 8'h00;
            15'd18392: data <= 8'h00;
            15'd18393: data <= 8'h00;
            15'd18394: data <= 8'h00;
            15'd18395: data <= 8'h03;
            15'd18396: data <= 8'hFF;
            15'd18397: data <= 8'hFE;
            15'd18398: data <= 8'h07;
            15'd18399: data <= 8'hFF;
            15'd18400: data <= 8'hFF;
            15'd18401: data <= 8'hFF;
            15'd18402: data <= 8'hFF;
            15'd18403: data <= 8'hFF;
            15'd18404: data <= 8'hFF;
            15'd18405: data <= 8'hFF;
            15'd18406: data <= 8'hFF;
            15'd18407: data <= 8'hFF;
            15'd18408: data <= 8'hFF;
            15'd18409: data <= 8'hFF;
            15'd18410: data <= 8'hFC;
            15'd18411: data <= 8'h07;
            15'd18412: data <= 8'hFF;
            15'd18413: data <= 8'hFF;
            15'd18414: data <= 8'h80;
            15'd18415: data <= 8'h00;
            15'd18416: data <= 8'h00;
            15'd18417: data <= 8'h00;
            15'd18418: data <= 8'h00;
            15'd18419: data <= 8'h00;
            15'd18420: data <= 8'h00;
            15'd18421: data <= 8'h00;
            15'd18422: data <= 8'h00;
            15'd18423: data <= 8'h00;
            15'd18424: data <= 8'h00;
            15'd18425: data <= 8'h03;
            15'd18426: data <= 8'hFF;
            15'd18427: data <= 8'hFE;
            15'd18428: data <= 8'h07;
            15'd18429: data <= 8'hFF;
            15'd18430: data <= 8'hFB;
            15'd18431: data <= 8'hFF;
            15'd18432: data <= 8'hFF;
            15'd18433: data <= 8'hFF;
            15'd18434: data <= 8'hFF;
            15'd18435: data <= 8'hFF;
            15'd18436: data <= 8'hFF;
            15'd18437: data <= 8'hFF;
            15'd18438: data <= 8'hFF;
            15'd18439: data <= 8'hFF;
            15'd18440: data <= 8'hFC;
            15'd18441: data <= 8'h07;
            15'd18442: data <= 8'hFF;
            15'd18443: data <= 8'hFF;
            15'd18444: data <= 8'h80;
            15'd18445: data <= 8'h00;
            15'd18446: data <= 8'h00;
            15'd18447: data <= 8'h00;
            15'd18448: data <= 8'h00;
            15'd18449: data <= 8'h00;
            15'd18450: data <= 8'h00;
            15'd18451: data <= 8'h00;
            15'd18452: data <= 8'h00;
            15'd18453: data <= 8'h00;
            15'd18454: data <= 8'h00;
            15'd18455: data <= 8'h03;
            15'd18456: data <= 8'hFF;
            15'd18457: data <= 8'hFF;
            15'd18458: data <= 8'h03;
            15'd18459: data <= 8'hFF;
            15'd18460: data <= 8'hF1;
            15'd18461: data <= 8'hFF;
            15'd18462: data <= 8'hFF;
            15'd18463: data <= 8'hFF;
            15'd18464: data <= 8'hFF;
            15'd18465: data <= 8'hFF;
            15'd18466: data <= 8'hFF;
            15'd18467: data <= 8'hFF;
            15'd18468: data <= 8'hFF;
            15'd18469: data <= 8'hFF;
            15'd18470: data <= 8'hFE;
            15'd18471: data <= 8'h03;
            15'd18472: data <= 8'hFF;
            15'd18473: data <= 8'hFF;
            15'd18474: data <= 8'h80;
            15'd18475: data <= 8'h00;
            15'd18476: data <= 8'h00;
            15'd18477: data <= 8'h00;
            15'd18478: data <= 8'h00;
            15'd18479: data <= 8'h00;
            15'd18480: data <= 8'h00;
            15'd18481: data <= 8'h00;
            15'd18482: data <= 8'h00;
            15'd18483: data <= 8'h00;
            15'd18484: data <= 8'h00;
            15'd18485: data <= 8'h03;
            15'd18486: data <= 8'hFF;
            15'd18487: data <= 8'hFF;
            15'd18488: data <= 8'h03;
            15'd18489: data <= 8'hFF;
            15'd18490: data <= 8'hE0;
            15'd18491: data <= 8'h38;
            15'd18492: data <= 8'h3F;
            15'd18493: data <= 8'hFF;
            15'd18494: data <= 8'hFF;
            15'd18495: data <= 8'hFF;
            15'd18496: data <= 8'hFF;
            15'd18497: data <= 8'hFF;
            15'd18498: data <= 8'hFF;
            15'd18499: data <= 8'hFF;
            15'd18500: data <= 8'hFE;
            15'd18501: data <= 8'h03;
            15'd18502: data <= 8'hFF;
            15'd18503: data <= 8'hFF;
            15'd18504: data <= 8'h80;
            15'd18505: data <= 8'h00;
            15'd18506: data <= 8'h00;
            15'd18507: data <= 8'h00;
            15'd18508: data <= 8'h00;
            15'd18509: data <= 8'h00;
            15'd18510: data <= 8'h00;
            15'd18511: data <= 8'h00;
            15'd18512: data <= 8'h00;
            15'd18513: data <= 8'h00;
            15'd18514: data <= 8'h00;
            15'd18515: data <= 8'h03;
            15'd18516: data <= 8'hFF;
            15'd18517: data <= 8'hFF;
            15'd18518: data <= 8'h83;
            15'd18519: data <= 8'hFF;
            15'd18520: data <= 8'hE0;
            15'd18521: data <= 8'h00;
            15'd18522: data <= 8'h3F;
            15'd18523: data <= 8'hFF;
            15'd18524: data <= 8'hFF;
            15'd18525: data <= 8'hFF;
            15'd18526: data <= 8'hFF;
            15'd18527: data <= 8'hFF;
            15'd18528: data <= 8'hFF;
            15'd18529: data <= 8'hFF;
            15'd18530: data <= 8'hFF;
            15'd18531: data <= 8'h01;
            15'd18532: data <= 8'hFF;
            15'd18533: data <= 8'hFF;
            15'd18534: data <= 8'h80;
            15'd18535: data <= 8'h00;
            15'd18536: data <= 8'h00;
            15'd18537: data <= 8'h00;
            15'd18538: data <= 8'h00;
            15'd18539: data <= 8'h00;
            15'd18540: data <= 8'h00;
            15'd18541: data <= 8'h00;
            15'd18542: data <= 8'h00;
            15'd18543: data <= 8'h00;
            15'd18544: data <= 8'h00;
            15'd18545: data <= 8'h03;
            15'd18546: data <= 8'hFF;
            15'd18547: data <= 8'hFF;
            15'd18548: data <= 8'h81;
            15'd18549: data <= 8'h03;
            15'd18550: data <= 8'hE0;
            15'd18551: data <= 8'h00;
            15'd18552: data <= 8'h3F;
            15'd18553: data <= 8'hFF;
            15'd18554: data <= 8'hFF;
            15'd18555: data <= 8'hFF;
            15'd18556: data <= 8'hFF;
            15'd18557: data <= 8'hFF;
            15'd18558: data <= 8'hFF;
            15'd18559: data <= 8'hFF;
            15'd18560: data <= 8'hFF;
            15'd18561: data <= 8'h00;
            15'd18562: data <= 8'hFF;
            15'd18563: data <= 8'hFF;
            15'd18564: data <= 8'h80;
            15'd18565: data <= 8'h00;
            15'd18566: data <= 8'h00;
            15'd18567: data <= 8'h00;
            15'd18568: data <= 8'h00;
            15'd18569: data <= 8'h00;
            15'd18570: data <= 8'h00;
            15'd18571: data <= 8'h00;
            15'd18572: data <= 8'h00;
            15'd18573: data <= 8'h00;
            15'd18574: data <= 8'h00;
            15'd18575: data <= 8'h03;
            15'd18576: data <= 8'hFF;
            15'd18577: data <= 8'hFF;
            15'd18578: data <= 8'hC0;
            15'd18579: data <= 8'h00;
            15'd18580: data <= 8'h70;
            15'd18581: data <= 8'h00;
            15'd18582: data <= 8'h1F;
            15'd18583: data <= 8'hFF;
            15'd18584: data <= 8'hFF;
            15'd18585: data <= 8'hFF;
            15'd18586: data <= 8'hFF;
            15'd18587: data <= 8'hFF;
            15'd18588: data <= 8'hFF;
            15'd18589: data <= 8'hFF;
            15'd18590: data <= 8'hFF;
            15'd18591: data <= 8'h80;
            15'd18592: data <= 8'h7F;
            15'd18593: data <= 8'hFF;
            15'd18594: data <= 8'h80;
            15'd18595: data <= 8'h00;
            15'd18596: data <= 8'h00;
            15'd18597: data <= 8'h00;
            15'd18598: data <= 8'h00;
            15'd18599: data <= 8'h00;
            15'd18600: data <= 8'h00;
            15'd18601: data <= 8'h00;
            15'd18602: data <= 8'h00;
            15'd18603: data <= 8'h00;
            15'd18604: data <= 8'h00;
            15'd18605: data <= 8'h03;
            15'd18606: data <= 8'hFF;
            15'd18607: data <= 8'hFF;
            15'd18608: data <= 8'hE0;
            15'd18609: data <= 8'h00;
            15'd18610: data <= 8'h18;
            15'd18611: data <= 8'h00;
            15'd18612: data <= 8'h7F;
            15'd18613: data <= 8'hFF;
            15'd18614: data <= 8'hFF;
            15'd18615: data <= 8'hFF;
            15'd18616: data <= 8'hFF;
            15'd18617: data <= 8'hFF;
            15'd18618: data <= 8'hFF;
            15'd18619: data <= 8'hFF;
            15'd18620: data <= 8'hFF;
            15'd18621: data <= 8'h80;
            15'd18622: data <= 8'h7F;
            15'd18623: data <= 8'hFF;
            15'd18624: data <= 8'h80;
            15'd18625: data <= 8'h00;
            15'd18626: data <= 8'h00;
            15'd18627: data <= 8'h00;
            15'd18628: data <= 8'h00;
            15'd18629: data <= 8'h00;
            15'd18630: data <= 8'h00;
            15'd18631: data <= 8'h00;
            15'd18632: data <= 8'h00;
            15'd18633: data <= 8'h00;
            15'd18634: data <= 8'h00;
            15'd18635: data <= 8'h03;
            15'd18636: data <= 8'hFF;
            15'd18637: data <= 8'hFF;
            15'd18638: data <= 8'hC0;
            15'd18639: data <= 8'h00;
            15'd18640: data <= 8'h03;
            15'd18641: data <= 8'hF3;
            15'd18642: data <= 8'hFF;
            15'd18643: data <= 8'hFF;
            15'd18644: data <= 8'hFF;
            15'd18645: data <= 8'hFF;
            15'd18646: data <= 8'hFF;
            15'd18647: data <= 8'hFF;
            15'd18648: data <= 8'hFF;
            15'd18649: data <= 8'hFF;
            15'd18650: data <= 8'hFF;
            15'd18651: data <= 8'hC0;
            15'd18652: data <= 8'h7F;
            15'd18653: data <= 8'hFF;
            15'd18654: data <= 8'h80;
            15'd18655: data <= 8'h00;
            15'd18656: data <= 8'h00;
            15'd18657: data <= 8'h00;
            15'd18658: data <= 8'h00;
            15'd18659: data <= 8'h00;
            15'd18660: data <= 8'h00;
            15'd18661: data <= 8'h00;
            15'd18662: data <= 8'h00;
            15'd18663: data <= 8'h00;
            15'd18664: data <= 8'h00;
            15'd18665: data <= 8'h03;
            15'd18666: data <= 8'hFF;
            15'd18667: data <= 8'hFF;
            15'd18668: data <= 8'hC0;
            15'd18669: data <= 8'h00;
            15'd18670: data <= 8'h01;
            15'd18671: data <= 8'hFF;
            15'd18672: data <= 8'hF8;
            15'd18673: data <= 8'h7F;
            15'd18674: data <= 8'hFF;
            15'd18675: data <= 8'hFF;
            15'd18676: data <= 8'hFF;
            15'd18677: data <= 8'hFF;
            15'd18678: data <= 8'hFF;
            15'd18679: data <= 8'hFF;
            15'd18680: data <= 8'hFF;
            15'd18681: data <= 8'hC0;
            15'd18682: data <= 8'h3F;
            15'd18683: data <= 8'hFF;
            15'd18684: data <= 8'h80;
            15'd18685: data <= 8'h00;
            15'd18686: data <= 8'h00;
            15'd18687: data <= 8'h00;
            15'd18688: data <= 8'h00;
            15'd18689: data <= 8'h00;
            15'd18690: data <= 8'h00;
            15'd18691: data <= 8'h00;
            15'd18692: data <= 8'h00;
            15'd18693: data <= 8'h00;
            15'd18694: data <= 8'h00;
            15'd18695: data <= 8'h03;
            15'd18696: data <= 8'hFF;
            15'd18697: data <= 8'hFF;
            15'd18698: data <= 8'hF0;
            15'd18699: data <= 8'h00;
            15'd18700: data <= 8'h00;
            15'd18701: data <= 8'h0F;
            15'd18702: data <= 8'hC0;
            15'd18703: data <= 8'h7F;
            15'd18704: data <= 8'hFF;
            15'd18705: data <= 8'hFF;
            15'd18706: data <= 8'hFF;
            15'd18707: data <= 8'hFF;
            15'd18708: data <= 8'hFF;
            15'd18709: data <= 8'hFF;
            15'd18710: data <= 8'hFF;
            15'd18711: data <= 8'hE0;
            15'd18712: data <= 8'h3F;
            15'd18713: data <= 8'hFF;
            15'd18714: data <= 8'h80;
            15'd18715: data <= 8'h00;
            15'd18716: data <= 8'h00;
            15'd18717: data <= 8'h00;
            15'd18718: data <= 8'h00;
            15'd18719: data <= 8'h00;
            15'd18720: data <= 8'h00;
            15'd18721: data <= 8'h00;
            15'd18722: data <= 8'h00;
            15'd18723: data <= 8'h00;
            15'd18724: data <= 8'h00;
            15'd18725: data <= 8'h03;
            15'd18726: data <= 8'hFF;
            15'd18727: data <= 8'hFF;
            15'd18728: data <= 8'hF8;
            15'd18729: data <= 8'h00;
            15'd18730: data <= 8'h00;
            15'd18731: data <= 8'h04;
            15'd18732: data <= 8'h00;
            15'd18733: data <= 8'h7F;
            15'd18734: data <= 8'hFF;
            15'd18735: data <= 8'hFF;
            15'd18736: data <= 8'hFF;
            15'd18737: data <= 8'hFF;
            15'd18738: data <= 8'hFF;
            15'd18739: data <= 8'hFF;
            15'd18740: data <= 8'hFF;
            15'd18741: data <= 8'hE0;
            15'd18742: data <= 8'h1F;
            15'd18743: data <= 8'hFF;
            15'd18744: data <= 8'h80;
            15'd18745: data <= 8'h00;
            15'd18746: data <= 8'h00;
            15'd18747: data <= 8'h00;
            15'd18748: data <= 8'h00;
            15'd18749: data <= 8'h00;
            15'd18750: data <= 8'h00;
            15'd18751: data <= 8'h00;
            15'd18752: data <= 8'h00;
            15'd18753: data <= 8'h00;
            15'd18754: data <= 8'h00;
            15'd18755: data <= 8'h03;
            15'd18756: data <= 8'hFF;
            15'd18757: data <= 8'hFF;
            15'd18758: data <= 8'hF8;
            15'd18759: data <= 8'h00;
            15'd18760: data <= 8'h00;
            15'd18761: data <= 8'h00;
            15'd18762: data <= 8'h00;
            15'd18763: data <= 8'hFF;
            15'd18764: data <= 8'hFF;
            15'd18765: data <= 8'hFF;
            15'd18766: data <= 8'hFF;
            15'd18767: data <= 8'hFF;
            15'd18768: data <= 8'hFF;
            15'd18769: data <= 8'hFF;
            15'd18770: data <= 8'hFF;
            15'd18771: data <= 8'hF0;
            15'd18772: data <= 8'h1F;
            15'd18773: data <= 8'hFF;
            15'd18774: data <= 8'h80;
            15'd18775: data <= 8'h00;
            15'd18776: data <= 8'h00;
            15'd18777: data <= 8'h00;
            15'd18778: data <= 8'h00;
            15'd18779: data <= 8'h00;
            15'd18780: data <= 8'h00;
            15'd18781: data <= 8'h00;
            15'd18782: data <= 8'h00;
            15'd18783: data <= 8'h00;
            15'd18784: data <= 8'h00;
            15'd18785: data <= 8'h03;
            15'd18786: data <= 8'hFF;
            15'd18787: data <= 8'hFF;
            15'd18788: data <= 8'hFE;
            15'd18789: data <= 8'h00;
            15'd18790: data <= 8'h08;
            15'd18791: data <= 8'h00;
            15'd18792: data <= 8'h01;
            15'd18793: data <= 8'hFF;
            15'd18794: data <= 8'hFF;
            15'd18795: data <= 8'hFF;
            15'd18796: data <= 8'hFF;
            15'd18797: data <= 8'hFF;
            15'd18798: data <= 8'hFF;
            15'd18799: data <= 8'hFF;
            15'd18800: data <= 8'hFF;
            15'd18801: data <= 8'hF0;
            15'd18802: data <= 8'h1F;
            15'd18803: data <= 8'hFF;
            15'd18804: data <= 8'h80;
            15'd18805: data <= 8'h00;
            15'd18806: data <= 8'h00;
            15'd18807: data <= 8'h00;
            15'd18808: data <= 8'h00;
            15'd18809: data <= 8'h00;
            15'd18810: data <= 8'h00;
            15'd18811: data <= 8'h00;
            15'd18812: data <= 8'h00;
            15'd18813: data <= 8'h00;
            15'd18814: data <= 8'h00;
            15'd18815: data <= 8'h03;
            15'd18816: data <= 8'hFF;
            15'd18817: data <= 8'hFF;
            15'd18818: data <= 8'hFF;
            15'd18819: data <= 8'h00;
            15'd18820: data <= 8'h04;
            15'd18821: data <= 8'h00;
            15'd18822: data <= 8'h01;
            15'd18823: data <= 8'hFF;
            15'd18824: data <= 8'hFF;
            15'd18825: data <= 8'hFF;
            15'd18826: data <= 8'hFF;
            15'd18827: data <= 8'hFF;
            15'd18828: data <= 8'hFF;
            15'd18829: data <= 8'hFF;
            15'd18830: data <= 8'hFF;
            15'd18831: data <= 8'hF8;
            15'd18832: data <= 8'h0F;
            15'd18833: data <= 8'hFF;
            15'd18834: data <= 8'h80;
            15'd18835: data <= 8'h00;
            15'd18836: data <= 8'h00;
            15'd18837: data <= 8'h00;
            15'd18838: data <= 8'h00;
            15'd18839: data <= 8'h00;
            15'd18840: data <= 8'h00;
            15'd18841: data <= 8'h00;
            15'd18842: data <= 8'h00;
            15'd18843: data <= 8'h00;
            15'd18844: data <= 8'h00;
            15'd18845: data <= 8'h03;
            15'd18846: data <= 8'hFF;
            15'd18847: data <= 8'hFF;
            15'd18848: data <= 8'hFF;
            15'd18849: data <= 8'h80;
            15'd18850: data <= 8'h07;
            15'd18851: data <= 8'h80;
            15'd18852: data <= 8'h03;
            15'd18853: data <= 8'hFF;
            15'd18854: data <= 8'hFF;
            15'd18855: data <= 8'hFF;
            15'd18856: data <= 8'hFF;
            15'd18857: data <= 8'hFF;
            15'd18858: data <= 8'hFF;
            15'd18859: data <= 8'hFF;
            15'd18860: data <= 8'hFF;
            15'd18861: data <= 8'hF8;
            15'd18862: data <= 8'h0F;
            15'd18863: data <= 8'hFF;
            15'd18864: data <= 8'h80;
            15'd18865: data <= 8'h00;
            15'd18866: data <= 8'h00;
            15'd18867: data <= 8'h00;
            15'd18868: data <= 8'h00;
            15'd18869: data <= 8'h00;
            15'd18870: data <= 8'h00;
            15'd18871: data <= 8'h00;
            15'd18872: data <= 8'h00;
            15'd18873: data <= 8'h00;
            15'd18874: data <= 8'h00;
            15'd18875: data <= 8'h03;
            15'd18876: data <= 8'hFF;
            15'd18877: data <= 8'hFF;
            15'd18878: data <= 8'hFF;
            15'd18879: data <= 8'hE0;
            15'd18880: data <= 8'h07;
            15'd18881: data <= 8'hFF;
            15'd18882: data <= 8'hC7;
            15'd18883: data <= 8'hFF;
            15'd18884: data <= 8'hFF;
            15'd18885: data <= 8'hFF;
            15'd18886: data <= 8'hFF;
            15'd18887: data <= 8'hFF;
            15'd18888: data <= 8'hFF;
            15'd18889: data <= 8'hFF;
            15'd18890: data <= 8'hFF;
            15'd18891: data <= 8'hFC;
            15'd18892: data <= 8'h07;
            15'd18893: data <= 8'hFF;
            15'd18894: data <= 8'h80;
            15'd18895: data <= 8'h00;
            15'd18896: data <= 8'h00;
            15'd18897: data <= 8'h00;
            15'd18898: data <= 8'h00;
            15'd18899: data <= 8'h00;
            15'd18900: data <= 8'h00;
            15'd18901: data <= 8'h00;
            15'd18902: data <= 8'h00;
            15'd18903: data <= 8'h00;
            15'd18904: data <= 8'h00;
            15'd18905: data <= 8'h03;
            15'd18906: data <= 8'hFF;
            15'd18907: data <= 8'hFF;
            15'd18908: data <= 8'hFF;
            15'd18909: data <= 8'hF0;
            15'd18910: data <= 8'h83;
            15'd18911: data <= 8'hFF;
            15'd18912: data <= 8'hC7;
            15'd18913: data <= 8'hFF;
            15'd18914: data <= 8'hFF;
            15'd18915: data <= 8'hFF;
            15'd18916: data <= 8'hFF;
            15'd18917: data <= 8'hFF;
            15'd18918: data <= 8'hFF;
            15'd18919: data <= 8'hFF;
            15'd18920: data <= 8'hFF;
            15'd18921: data <= 8'hFC;
            15'd18922: data <= 8'h07;
            15'd18923: data <= 8'hFF;
            15'd18924: data <= 8'h80;
            15'd18925: data <= 8'h00;
            15'd18926: data <= 8'h00;
            15'd18927: data <= 8'h00;
            15'd18928: data <= 8'h00;
            15'd18929: data <= 8'h00;
            15'd18930: data <= 8'h00;
            15'd18931: data <= 8'h00;
            15'd18932: data <= 8'h00;
            15'd18933: data <= 8'h00;
            15'd18934: data <= 8'h00;
            15'd18935: data <= 8'h03;
            15'd18936: data <= 8'hFF;
            15'd18937: data <= 8'hFF;
            15'd18938: data <= 8'hFF;
            15'd18939: data <= 8'hF0;
            15'd18940: data <= 8'hC1;
            15'd18941: data <= 8'hFF;
            15'd18942: data <= 8'hC7;
            15'd18943: data <= 8'hFF;
            15'd18944: data <= 8'hFF;
            15'd18945: data <= 8'hFF;
            15'd18946: data <= 8'hFF;
            15'd18947: data <= 8'hFF;
            15'd18948: data <= 8'hFF;
            15'd18949: data <= 8'hFF;
            15'd18950: data <= 8'hFF;
            15'd18951: data <= 8'hFC;
            15'd18952: data <= 8'h07;
            15'd18953: data <= 8'hFF;
            15'd18954: data <= 8'h80;
            15'd18955: data <= 8'h00;
            15'd18956: data <= 8'h00;
            15'd18957: data <= 8'h00;
            15'd18958: data <= 8'h00;
            15'd18959: data <= 8'h00;
            15'd18960: data <= 8'h00;
            15'd18961: data <= 8'h00;
            15'd18962: data <= 8'h00;
            15'd18963: data <= 8'h00;
            15'd18964: data <= 8'h00;
            15'd18965: data <= 8'h03;
            15'd18966: data <= 8'hFF;
            15'd18967: data <= 8'hFF;
            15'd18968: data <= 8'hFF;
            15'd18969: data <= 8'hF0;
            15'd18970: data <= 8'hE1;
            15'd18971: data <= 8'hFF;
            15'd18972: data <= 8'hC7;
            15'd18973: data <= 8'hFF;
            15'd18974: data <= 8'hFF;
            15'd18975: data <= 8'hFF;
            15'd18976: data <= 8'hFF;
            15'd18977: data <= 8'hFF;
            15'd18978: data <= 8'hFF;
            15'd18979: data <= 8'hFF;
            15'd18980: data <= 8'hFF;
            15'd18981: data <= 8'hFE;
            15'd18982: data <= 8'h03;
            15'd18983: data <= 8'hFF;
            15'd18984: data <= 8'h80;
            15'd18985: data <= 8'h00;
            15'd18986: data <= 8'h00;
            15'd18987: data <= 8'h00;
            15'd18988: data <= 8'h00;
            15'd18989: data <= 8'h00;
            15'd18990: data <= 8'h00;
            15'd18991: data <= 8'h00;
            15'd18992: data <= 8'h00;
            15'd18993: data <= 8'h00;
            15'd18994: data <= 8'h00;
            15'd18995: data <= 8'h03;
            15'd18996: data <= 8'hFF;
            15'd18997: data <= 8'hFF;
            15'd18998: data <= 8'hFF;
            15'd18999: data <= 8'hF0;
            15'd19000: data <= 8'hF0;
            15'd19001: data <= 8'hFF;
            15'd19002: data <= 8'hC7;
            15'd19003: data <= 8'hFF;
            15'd19004: data <= 8'hFF;
            15'd19005: data <= 8'hFF;
            15'd19006: data <= 8'hFF;
            15'd19007: data <= 8'hFF;
            15'd19008: data <= 8'hFF;
            15'd19009: data <= 8'hFF;
            15'd19010: data <= 8'hFF;
            15'd19011: data <= 8'hFE;
            15'd19012: data <= 8'h03;
            15'd19013: data <= 8'hFF;
            15'd19014: data <= 8'h80;
            15'd19015: data <= 8'h00;
            15'd19016: data <= 8'h00;
            15'd19017: data <= 8'h00;
            15'd19018: data <= 8'h00;
            15'd19019: data <= 8'h00;
            15'd19020: data <= 8'h00;
            15'd19021: data <= 8'h00;
            15'd19022: data <= 8'h00;
            15'd19023: data <= 8'h00;
            15'd19024: data <= 8'h00;
            15'd19025: data <= 8'h03;
            15'd19026: data <= 8'hFF;
            15'd19027: data <= 8'hFF;
            15'd19028: data <= 8'hFF;
            15'd19029: data <= 8'hF8;
            15'd19030: data <= 8'h70;
            15'd19031: data <= 8'hFF;
            15'd19032: data <= 8'hE3;
            15'd19033: data <= 8'hFF;
            15'd19034: data <= 8'hFF;
            15'd19035: data <= 8'hFF;
            15'd19036: data <= 8'hFF;
            15'd19037: data <= 8'hFF;
            15'd19038: data <= 8'hFF;
            15'd19039: data <= 8'hFF;
            15'd19040: data <= 8'hFF;
            15'd19041: data <= 8'hFF;
            15'd19042: data <= 8'h01;
            15'd19043: data <= 8'hFF;
            15'd19044: data <= 8'h80;
            15'd19045: data <= 8'h00;
            15'd19046: data <= 8'h00;
            15'd19047: data <= 8'h00;
            15'd19048: data <= 8'h00;
            15'd19049: data <= 8'h00;
            15'd19050: data <= 8'h00;
            15'd19051: data <= 8'h00;
            15'd19052: data <= 8'h00;
            15'd19053: data <= 8'h00;
            15'd19054: data <= 8'h00;
            15'd19055: data <= 8'h03;
            15'd19056: data <= 8'hFF;
            15'd19057: data <= 8'hFF;
            15'd19058: data <= 8'hFF;
            15'd19059: data <= 8'hF0;
            15'd19060: data <= 8'h78;
            15'd19061: data <= 8'hFF;
            15'd19062: data <= 8'hE1;
            15'd19063: data <= 8'hFF;
            15'd19064: data <= 8'hFF;
            15'd19065: data <= 8'hFF;
            15'd19066: data <= 8'hFF;
            15'd19067: data <= 8'hFF;
            15'd19068: data <= 8'hFF;
            15'd19069: data <= 8'hFF;
            15'd19070: data <= 8'hFF;
            15'd19071: data <= 8'hFF;
            15'd19072: data <= 8'h01;
            15'd19073: data <= 8'hFF;
            15'd19074: data <= 8'h80;
            15'd19075: data <= 8'h00;
            15'd19076: data <= 8'h00;
            15'd19077: data <= 8'h00;
            15'd19078: data <= 8'h00;
            15'd19079: data <= 8'h00;
            15'd19080: data <= 8'h00;
            15'd19081: data <= 8'h00;
            15'd19082: data <= 8'h00;
            15'd19083: data <= 8'h00;
            15'd19084: data <= 8'h00;
            15'd19085: data <= 8'h03;
            15'd19086: data <= 8'hFF;
            15'd19087: data <= 8'hFF;
            15'd19088: data <= 8'hFF;
            15'd19089: data <= 8'hF0;
            15'd19090: data <= 8'h78;
            15'd19091: data <= 8'h7F;
            15'd19092: data <= 8'hE0;
            15'd19093: data <= 8'hFF;
            15'd19094: data <= 8'hFF;
            15'd19095: data <= 8'hFF;
            15'd19096: data <= 8'hFF;
            15'd19097: data <= 8'hFF;
            15'd19098: data <= 8'hFF;
            15'd19099: data <= 8'hFF;
            15'd19100: data <= 8'hFF;
            15'd19101: data <= 8'hFF;
            15'd19102: data <= 8'h80;
            15'd19103: data <= 8'hFF;
            15'd19104: data <= 8'h80;
            15'd19105: data <= 8'h00;
            15'd19106: data <= 8'h00;
            15'd19107: data <= 8'h00;
            15'd19108: data <= 8'h00;
            15'd19109: data <= 8'h00;
            15'd19110: data <= 8'h00;
            15'd19111: data <= 8'h00;
            15'd19112: data <= 8'h00;
            15'd19113: data <= 8'h00;
            15'd19114: data <= 8'h00;
            15'd19115: data <= 8'h03;
            15'd19116: data <= 8'hFF;
            15'd19117: data <= 8'hFF;
            15'd19118: data <= 8'hFF;
            15'd19119: data <= 8'hF0;
            15'd19120: data <= 8'h78;
            15'd19121: data <= 8'h7F;
            15'd19122: data <= 8'hE0;
            15'd19123: data <= 8'h7F;
            15'd19124: data <= 8'hFF;
            15'd19125: data <= 8'hFF;
            15'd19126: data <= 8'hFF;
            15'd19127: data <= 8'hFF;
            15'd19128: data <= 8'hFF;
            15'd19129: data <= 8'hFF;
            15'd19130: data <= 8'hFF;
            15'd19131: data <= 8'hFF;
            15'd19132: data <= 8'h80;
            15'd19133: data <= 8'hFF;
            15'd19134: data <= 8'h80;
            15'd19135: data <= 8'h00;
            15'd19136: data <= 8'h00;
            15'd19137: data <= 8'h00;
            15'd19138: data <= 8'h00;
            15'd19139: data <= 8'h00;
            15'd19140: data <= 8'h00;
            15'd19141: data <= 8'h00;
            15'd19142: data <= 8'h00;
            15'd19143: data <= 8'h00;
            15'd19144: data <= 8'h00;
            15'd19145: data <= 8'h03;
            15'd19146: data <= 8'hFF;
            15'd19147: data <= 8'hFF;
            15'd19148: data <= 8'hFF;
            15'd19149: data <= 8'hF0;
            15'd19150: data <= 8'h7C;
            15'd19151: data <= 8'h3F;
            15'd19152: data <= 8'hF0;
            15'd19153: data <= 8'h3F;
            15'd19154: data <= 8'hFF;
            15'd19155: data <= 8'hFF;
            15'd19156: data <= 8'hF0;
            15'd19157: data <= 8'h7F;
            15'd19158: data <= 8'hFF;
            15'd19159: data <= 8'hFF;
            15'd19160: data <= 8'hFF;
            15'd19161: data <= 8'hFF;
            15'd19162: data <= 8'hC0;
            15'd19163: data <= 8'h7F;
            15'd19164: data <= 8'h80;
            15'd19165: data <= 8'h00;
            15'd19166: data <= 8'h00;
            15'd19167: data <= 8'h00;
            15'd19168: data <= 8'h00;
            15'd19169: data <= 8'h00;
            15'd19170: data <= 8'h00;
            15'd19171: data <= 8'h00;
            15'd19172: data <= 8'h00;
            15'd19173: data <= 8'h00;
            15'd19174: data <= 8'h00;
            15'd19175: data <= 8'h03;
            15'd19176: data <= 8'hFF;
            15'd19177: data <= 8'hFF;
            15'd19178: data <= 8'hFF;
            15'd19179: data <= 8'hF8;
            15'd19180: data <= 8'h7C;
            15'd19181: data <= 8'h3F;
            15'd19182: data <= 8'hF8;
            15'd19183: data <= 8'h0F;
            15'd19184: data <= 8'hFF;
            15'd19185: data <= 8'hFF;
            15'd19186: data <= 8'hE0;
            15'd19187: data <= 8'h7F;
            15'd19188: data <= 8'hFF;
            15'd19189: data <= 8'hFF;
            15'd19190: data <= 8'hFF;
            15'd19191: data <= 8'hFF;
            15'd19192: data <= 8'hC0;
            15'd19193: data <= 8'h7F;
            15'd19194: data <= 8'h80;
            15'd19195: data <= 8'h00;
            15'd19196: data <= 8'h00;
            15'd19197: data <= 8'h00;
            15'd19198: data <= 8'h00;
            15'd19199: data <= 8'h00;
            15'd19200: data <= 8'h00;
            15'd19201: data <= 8'h00;
            15'd19202: data <= 8'h00;
            15'd19203: data <= 8'h00;
            15'd19204: data <= 8'h00;
            15'd19205: data <= 8'h03;
            15'd19206: data <= 8'hFF;
            15'd19207: data <= 8'hFF;
            15'd19208: data <= 8'hFF;
            15'd19209: data <= 8'hF8;
            15'd19210: data <= 8'h7C;
            15'd19211: data <= 8'h3F;
            15'd19212: data <= 8'hFC;
            15'd19213: data <= 8'h03;
            15'd19214: data <= 8'hFF;
            15'd19215: data <= 8'hFF;
            15'd19216: data <= 8'hC0;
            15'd19217: data <= 8'h7F;
            15'd19218: data <= 8'hFF;
            15'd19219: data <= 8'hFF;
            15'd19220: data <= 8'hFF;
            15'd19221: data <= 8'hFF;
            15'd19222: data <= 8'hC0;
            15'd19223: data <= 8'h7F;
            15'd19224: data <= 8'h80;
            15'd19225: data <= 8'h00;
            15'd19226: data <= 8'h00;
            15'd19227: data <= 8'h00;
            15'd19228: data <= 8'h00;
            15'd19229: data <= 8'h00;
            15'd19230: data <= 8'h00;
            15'd19231: data <= 8'h00;
            15'd19232: data <= 8'h00;
            15'd19233: data <= 8'h00;
            15'd19234: data <= 8'h00;
            15'd19235: data <= 8'h03;
            15'd19236: data <= 8'hFF;
            15'd19237: data <= 8'hFF;
            15'd19238: data <= 8'hFF;
            15'd19239: data <= 8'hFC;
            15'd19240: data <= 8'h7C;
            15'd19241: data <= 8'h3F;
            15'd19242: data <= 8'hFE;
            15'd19243: data <= 8'h00;
            15'd19244: data <= 8'hFF;
            15'd19245: data <= 8'hFF;
            15'd19246: data <= 8'h00;
            15'd19247: data <= 8'h7F;
            15'd19248: data <= 8'hFF;
            15'd19249: data <= 8'hFF;
            15'd19250: data <= 8'hFF;
            15'd19251: data <= 8'hFF;
            15'd19252: data <= 8'hE0;
            15'd19253: data <= 8'h3F;
            15'd19254: data <= 8'h80;
            15'd19255: data <= 8'h00;
            15'd19256: data <= 8'h00;
            15'd19257: data <= 8'h00;
            15'd19258: data <= 8'h00;
            15'd19259: data <= 8'h00;
            15'd19260: data <= 8'h00;
            15'd19261: data <= 8'h00;
            15'd19262: data <= 8'h00;
            15'd19263: data <= 8'h00;
            15'd19264: data <= 8'h00;
            15'd19265: data <= 8'h03;
            15'd19266: data <= 8'hFF;
            15'd19267: data <= 8'hFF;
            15'd19268: data <= 8'hFF;
            15'd19269: data <= 8'hFC;
            15'd19270: data <= 8'h7C;
            15'd19271: data <= 8'h1F;
            15'd19272: data <= 8'hFF;
            15'd19273: data <= 8'h80;
            15'd19274: data <= 8'h1F;
            15'd19275: data <= 8'hFE;
            15'd19276: data <= 8'h00;
            15'd19277: data <= 8'h7F;
            15'd19278: data <= 8'hFF;
            15'd19279: data <= 8'hFF;
            15'd19280: data <= 8'hFF;
            15'd19281: data <= 8'hFF;
            15'd19282: data <= 8'hE0;
            15'd19283: data <= 8'h3F;
            15'd19284: data <= 8'h80;
            15'd19285: data <= 8'h00;
            15'd19286: data <= 8'h00;
            15'd19287: data <= 8'h00;
            15'd19288: data <= 8'h00;
            15'd19289: data <= 8'h00;
            15'd19290: data <= 8'h00;
            15'd19291: data <= 8'h00;
            15'd19292: data <= 8'h00;
            15'd19293: data <= 8'h00;
            15'd19294: data <= 8'h00;
            15'd19295: data <= 8'h03;
            15'd19296: data <= 8'hFF;
            15'd19297: data <= 8'hFF;
            15'd19298: data <= 8'hFF;
            15'd19299: data <= 8'hF8;
            15'd19300: data <= 8'h7E;
            15'd19301: data <= 8'h1F;
            15'd19302: data <= 8'hFF;
            15'd19303: data <= 8'hC0;
            15'd19304: data <= 8'h03;
            15'd19305: data <= 8'h00;
            15'd19306: data <= 8'h00;
            15'd19307: data <= 8'hFF;
            15'd19308: data <= 8'hFF;
            15'd19309: data <= 8'hFF;
            15'd19310: data <= 8'hFF;
            15'd19311: data <= 8'hFF;
            15'd19312: data <= 8'hE0;
            15'd19313: data <= 8'h1F;
            15'd19314: data <= 8'h80;
            15'd19315: data <= 8'h00;
            15'd19316: data <= 8'h00;
            15'd19317: data <= 8'h00;
            15'd19318: data <= 8'h00;
            15'd19319: data <= 8'h00;
            15'd19320: data <= 8'h00;
            15'd19321: data <= 8'h00;
            15'd19322: data <= 8'h00;
            15'd19323: data <= 8'h00;
            15'd19324: data <= 8'h00;
            15'd19325: data <= 8'h03;
            15'd19326: data <= 8'hFF;
            15'd19327: data <= 8'hFF;
            15'd19328: data <= 8'hFF;
            15'd19329: data <= 8'hF8;
            15'd19330: data <= 8'h7E;
            15'd19331: data <= 8'h0F;
            15'd19332: data <= 8'hFF;
            15'd19333: data <= 8'hE0;
            15'd19334: data <= 8'h00;
            15'd19335: data <= 8'h00;
            15'd19336: data <= 8'h03;
            15'd19337: data <= 8'hFF;
            15'd19338: data <= 8'hFF;
            15'd19339: data <= 8'hFF;
            15'd19340: data <= 8'hFF;
            15'd19341: data <= 8'hFF;
            15'd19342: data <= 8'hE0;
            15'd19343: data <= 8'h1F;
            15'd19344: data <= 8'h80;
            15'd19345: data <= 8'h00;
            15'd19346: data <= 8'h00;
            15'd19347: data <= 8'h00;
            15'd19348: data <= 8'h00;
            15'd19349: data <= 8'h00;
            15'd19350: data <= 8'h00;
            15'd19351: data <= 8'h00;
            15'd19352: data <= 8'h00;
            15'd19353: data <= 8'h00;
            15'd19354: data <= 8'h00;
            15'd19355: data <= 8'h03;
            15'd19356: data <= 8'hFF;
            15'd19357: data <= 8'hFF;
            15'd19358: data <= 8'hFF;
            15'd19359: data <= 8'hF8;
            15'd19360: data <= 8'h7F;
            15'd19361: data <= 8'h0F;
            15'd19362: data <= 8'hFF;
            15'd19363: data <= 8'hF8;
            15'd19364: data <= 8'h00;
            15'd19365: data <= 8'h00;
            15'd19366: data <= 8'h07;
            15'd19367: data <= 8'hFF;
            15'd19368: data <= 8'hFF;
            15'd19369: data <= 8'hFF;
            15'd19370: data <= 8'hFF;
            15'd19371: data <= 8'hFF;
            15'd19372: data <= 8'hF0;
            15'd19373: data <= 8'h1F;
            15'd19374: data <= 8'h80;
            15'd19375: data <= 8'h00;
            15'd19376: data <= 8'h00;
            15'd19377: data <= 8'h00;
            15'd19378: data <= 8'h00;
            15'd19379: data <= 8'h00;
            15'd19380: data <= 8'h00;
            15'd19381: data <= 8'h00;
            15'd19382: data <= 8'h00;
            15'd19383: data <= 8'h00;
            15'd19384: data <= 8'h00;
            15'd19385: data <= 8'h03;
            15'd19386: data <= 8'hFF;
            15'd19387: data <= 8'hFF;
            15'd19388: data <= 8'hFF;
            15'd19389: data <= 8'hF8;
            15'd19390: data <= 8'h7F;
            15'd19391: data <= 8'h07;
            15'd19392: data <= 8'hFF;
            15'd19393: data <= 8'hFF;
            15'd19394: data <= 8'h00;
            15'd19395: data <= 8'h00;
            15'd19396: data <= 8'h1F;
            15'd19397: data <= 8'hFF;
            15'd19398: data <= 8'hFF;
            15'd19399: data <= 8'hFF;
            15'd19400: data <= 8'hFF;
            15'd19401: data <= 8'hFF;
            15'd19402: data <= 8'hF0;
            15'd19403: data <= 8'h1F;
            15'd19404: data <= 8'h80;
            15'd19405: data <= 8'h00;
            15'd19406: data <= 8'h00;
            15'd19407: data <= 8'h00;
            15'd19408: data <= 8'h00;
            15'd19409: data <= 8'h00;
            15'd19410: data <= 8'h00;
            15'd19411: data <= 8'h00;
            15'd19412: data <= 8'h00;
            15'd19413: data <= 8'h00;
            15'd19414: data <= 8'h00;
            15'd19415: data <= 8'h03;
            15'd19416: data <= 8'hFF;
            15'd19417: data <= 8'hFF;
            15'd19418: data <= 8'hFF;
            15'd19419: data <= 8'hF8;
            15'd19420: data <= 8'h7F;
            15'd19421: data <= 8'h87;
            15'd19422: data <= 8'hFF;
            15'd19423: data <= 8'hFF;
            15'd19424: data <= 8'hF0;
            15'd19425: data <= 8'h00;
            15'd19426: data <= 8'h7F;
            15'd19427: data <= 8'hFF;
            15'd19428: data <= 8'hFF;
            15'd19429: data <= 8'hFF;
            15'd19430: data <= 8'hFF;
            15'd19431: data <= 8'hFF;
            15'd19432: data <= 8'hF8;
            15'd19433: data <= 8'h0F;
            15'd19434: data <= 8'h80;
            15'd19435: data <= 8'h00;
            15'd19436: data <= 8'h00;
            15'd19437: data <= 8'h00;
            15'd19438: data <= 8'h00;
            15'd19439: data <= 8'h00;
            15'd19440: data <= 8'h00;
            15'd19441: data <= 8'h00;
            15'd19442: data <= 8'h00;
            15'd19443: data <= 8'h00;
            15'd19444: data <= 8'h00;
            15'd19445: data <= 8'h03;
            15'd19446: data <= 8'hFF;
            15'd19447: data <= 8'hFF;
            15'd19448: data <= 8'hFF;
            15'd19449: data <= 8'hF8;
            15'd19450: data <= 8'h7F;
            15'd19451: data <= 8'h83;
            15'd19452: data <= 8'hFF;
            15'd19453: data <= 8'hFF;
            15'd19454: data <= 8'hFE;
            15'd19455: data <= 8'h01;
            15'd19456: data <= 8'hFF;
            15'd19457: data <= 8'hFF;
            15'd19458: data <= 8'hFF;
            15'd19459: data <= 8'hFF;
            15'd19460: data <= 8'hFF;
            15'd19461: data <= 8'hFF;
            15'd19462: data <= 8'hF8;
            15'd19463: data <= 8'h0F;
            15'd19464: data <= 8'h80;
            15'd19465: data <= 8'h00;
            15'd19466: data <= 8'h00;
            15'd19467: data <= 8'h00;
            15'd19468: data <= 8'h00;
            15'd19469: data <= 8'h00;
            15'd19470: data <= 8'h00;
            15'd19471: data <= 8'h00;
            15'd19472: data <= 8'h00;
            15'd19473: data <= 8'h00;
            15'd19474: data <= 8'h00;
            15'd19475: data <= 8'h03;
            15'd19476: data <= 8'hFF;
            15'd19477: data <= 8'hFF;
            15'd19478: data <= 8'hFF;
            15'd19479: data <= 8'hF8;
            15'd19480: data <= 8'h7F;
            15'd19481: data <= 8'hC1;
            15'd19482: data <= 8'hFF;
            15'd19483: data <= 8'hFF;
            15'd19484: data <= 8'hFF;
            15'd19485: data <= 8'hFF;
            15'd19486: data <= 8'hFF;
            15'd19487: data <= 8'hFF;
            15'd19488: data <= 8'hFF;
            15'd19489: data <= 8'hFF;
            15'd19490: data <= 8'hFF;
            15'd19491: data <= 8'hFF;
            15'd19492: data <= 8'hF8;
            15'd19493: data <= 8'h0F;
            15'd19494: data <= 8'h80;
            15'd19495: data <= 8'h00;
            15'd19496: data <= 8'h00;
            15'd19497: data <= 8'h00;
            15'd19498: data <= 8'h00;
            15'd19499: data <= 8'h00;
            15'd19500: data <= 8'h00;
            15'd19501: data <= 8'h00;
            15'd19502: data <= 8'h00;
            15'd19503: data <= 8'h00;
            15'd19504: data <= 8'h00;
            15'd19505: data <= 8'h03;
            15'd19506: data <= 8'hFF;
            15'd19507: data <= 8'hFF;
            15'd19508: data <= 8'hFF;
            15'd19509: data <= 8'hF8;
            15'd19510: data <= 8'h7F;
            15'd19511: data <= 8'hC1;
            15'd19512: data <= 8'hFF;
            15'd19513: data <= 8'hFF;
            15'd19514: data <= 8'hFF;
            15'd19515: data <= 8'hFF;
            15'd19516: data <= 8'hFF;
            15'd19517: data <= 8'hFF;
            15'd19518: data <= 8'hFF;
            15'd19519: data <= 8'hFF;
            15'd19520: data <= 8'hFF;
            15'd19521: data <= 8'hFF;
            15'd19522: data <= 8'hF8;
            15'd19523: data <= 8'h07;
            15'd19524: data <= 8'h80;
            15'd19525: data <= 8'h00;
            15'd19526: data <= 8'h00;
            15'd19527: data <= 8'h00;
            15'd19528: data <= 8'h00;
            15'd19529: data <= 8'h00;
            15'd19530: data <= 8'h00;
            15'd19531: data <= 8'h00;
            15'd19532: data <= 8'h00;
            15'd19533: data <= 8'h00;
            15'd19534: data <= 8'h00;
            15'd19535: data <= 8'h03;
            15'd19536: data <= 8'hFF;
            15'd19537: data <= 8'hFF;
            15'd19538: data <= 8'hFF;
            15'd19539: data <= 8'hF8;
            15'd19540: data <= 8'h7F;
            15'd19541: data <= 8'hE0;
            15'd19542: data <= 8'hFF;
            15'd19543: data <= 8'hFF;
            15'd19544: data <= 8'hFF;
            15'd19545: data <= 8'hFF;
            15'd19546: data <= 8'hFF;
            15'd19547: data <= 8'hFF;
            15'd19548: data <= 8'hFF;
            15'd19549: data <= 8'hFF;
            15'd19550: data <= 8'hFF;
            15'd19551: data <= 8'hFF;
            15'd19552: data <= 8'hFC;
            15'd19553: data <= 8'h07;
            15'd19554: data <= 8'h80;
            15'd19555: data <= 8'h00;
            15'd19556: data <= 8'h00;
            15'd19557: data <= 8'h00;
            15'd19558: data <= 8'h00;
            15'd19559: data <= 8'h00;
            15'd19560: data <= 8'h00;
            15'd19561: data <= 8'h00;
            15'd19562: data <= 8'h00;
            15'd19563: data <= 8'h00;
            15'd19564: data <= 8'h00;
            15'd19565: data <= 8'h03;
            15'd19566: data <= 8'hFF;
            15'd19567: data <= 8'hFF;
            15'd19568: data <= 8'hFF;
            15'd19569: data <= 8'hFC;
            15'd19570: data <= 8'h7F;
            15'd19571: data <= 8'hE0;
            15'd19572: data <= 8'h7F;
            15'd19573: data <= 8'hFF;
            15'd19574: data <= 8'hFF;
            15'd19575: data <= 8'hFF;
            15'd19576: data <= 8'hFF;
            15'd19577: data <= 8'hFF;
            15'd19578: data <= 8'hFF;
            15'd19579: data <= 8'hFF;
            15'd19580: data <= 8'hFF;
            15'd19581: data <= 8'hFF;
            15'd19582: data <= 8'hFC;
            15'd19583: data <= 8'h07;
            15'd19584: data <= 8'h80;
            15'd19585: data <= 8'h00;
            15'd19586: data <= 8'h00;
            15'd19587: data <= 8'h00;
            15'd19588: data <= 8'h00;
            15'd19589: data <= 8'h00;
            15'd19590: data <= 8'h00;
            15'd19591: data <= 8'h00;
            15'd19592: data <= 8'h00;
            15'd19593: data <= 8'h00;
            15'd19594: data <= 8'h00;
            15'd19595: data <= 8'h03;
            15'd19596: data <= 8'hFF;
            15'd19597: data <= 8'hFF;
            15'd19598: data <= 8'hFF;
            15'd19599: data <= 8'hFC;
            15'd19600: data <= 8'h7F;
            15'd19601: data <= 8'hF0;
            15'd19602: data <= 8'h7F;
            15'd19603: data <= 8'hFF;
            15'd19604: data <= 8'hFF;
            15'd19605: data <= 8'hFF;
            15'd19606: data <= 8'hFF;
            15'd19607: data <= 8'hFF;
            15'd19608: data <= 8'hFF;
            15'd19609: data <= 8'hFF;
            15'd19610: data <= 8'hFF;
            15'd19611: data <= 8'hFF;
            15'd19612: data <= 8'hFC;
            15'd19613: data <= 8'h03;
            15'd19614: data <= 8'h80;
            15'd19615: data <= 8'h00;
            15'd19616: data <= 8'h00;
            15'd19617: data <= 8'h00;
            15'd19618: data <= 8'h00;
            15'd19619: data <= 8'h00;
            15'd19620: data <= 8'h00;
            15'd19621: data <= 8'h00;
            15'd19622: data <= 8'h00;
            15'd19623: data <= 8'h00;
            15'd19624: data <= 8'h00;
            15'd19625: data <= 8'h03;
            15'd19626: data <= 8'hFF;
            15'd19627: data <= 8'hFF;
            15'd19628: data <= 8'hFF;
            15'd19629: data <= 8'hFC;
            15'd19630: data <= 8'h7F;
            15'd19631: data <= 8'hF8;
            15'd19632: data <= 8'h3F;
            15'd19633: data <= 8'hFF;
            15'd19634: data <= 8'hFF;
            15'd19635: data <= 8'hFF;
            15'd19636: data <= 8'hFF;
            15'd19637: data <= 8'hFF;
            15'd19638: data <= 8'hFF;
            15'd19639: data <= 8'hFF;
            15'd19640: data <= 8'hFF;
            15'd19641: data <= 8'hFF;
            15'd19642: data <= 8'hFE;
            15'd19643: data <= 8'h03;
            15'd19644: data <= 8'h80;
            15'd19645: data <= 8'h00;
            15'd19646: data <= 8'h00;
            15'd19647: data <= 8'h00;
            15'd19648: data <= 8'h00;
            15'd19649: data <= 8'h00;
            15'd19650: data <= 8'h00;
            15'd19651: data <= 8'h00;
            15'd19652: data <= 8'h00;
            15'd19653: data <= 8'h00;
            15'd19654: data <= 8'h00;
            15'd19655: data <= 8'h03;
            15'd19656: data <= 8'hFF;
            15'd19657: data <= 8'hFF;
            15'd19658: data <= 8'hFF;
            15'd19659: data <= 8'hFC;
            15'd19660: data <= 8'h7F;
            15'd19661: data <= 8'hFC;
            15'd19662: data <= 8'h1F;
            15'd19663: data <= 8'hFF;
            15'd19664: data <= 8'hFF;
            15'd19665: data <= 8'hFF;
            15'd19666: data <= 8'hFF;
            15'd19667: data <= 8'hFF;
            15'd19668: data <= 8'hFF;
            15'd19669: data <= 8'hFF;
            15'd19670: data <= 8'hFF;
            15'd19671: data <= 8'hFF;
            15'd19672: data <= 8'hFE;
            15'd19673: data <= 8'h03;
            15'd19674: data <= 8'h80;
            15'd19675: data <= 8'h00;
            15'd19676: data <= 8'h00;
            15'd19677: data <= 8'h00;
            15'd19678: data <= 8'h00;
            15'd19679: data <= 8'h00;
            15'd19680: data <= 8'h00;
            15'd19681: data <= 8'h00;
            15'd19682: data <= 8'h00;
            15'd19683: data <= 8'h00;
            15'd19684: data <= 8'h00;
            15'd19685: data <= 8'h03;
            15'd19686: data <= 8'hFF;
            15'd19687: data <= 8'hFF;
            15'd19688: data <= 8'hFF;
            15'd19689: data <= 8'hFC;
            15'd19690: data <= 8'h7F;
            15'd19691: data <= 8'hFC;
            15'd19692: data <= 8'h0F;
            15'd19693: data <= 8'hFF;
            15'd19694: data <= 8'hFF;
            15'd19695: data <= 8'hFF;
            15'd19696: data <= 8'hFF;
            15'd19697: data <= 8'hFF;
            15'd19698: data <= 8'hFF;
            15'd19699: data <= 8'hFF;
            15'd19700: data <= 8'hFF;
            15'd19701: data <= 8'hFF;
            15'd19702: data <= 8'hFE;
            15'd19703: data <= 8'h03;
            15'd19704: data <= 8'h80;
            15'd19705: data <= 8'h00;
            15'd19706: data <= 8'h00;
            15'd19707: data <= 8'h00;
            15'd19708: data <= 8'h00;
            15'd19709: data <= 8'h00;
            15'd19710: data <= 8'h00;
            15'd19711: data <= 8'h00;
            15'd19712: data <= 8'h00;
            15'd19713: data <= 8'h00;
            15'd19714: data <= 8'h00;
            15'd19715: data <= 8'h03;
            15'd19716: data <= 8'hFF;
            15'd19717: data <= 8'hFF;
            15'd19718: data <= 8'hFF;
            15'd19719: data <= 8'hFC;
            15'd19720: data <= 8'h7F;
            15'd19721: data <= 8'hFE;
            15'd19722: data <= 8'h07;
            15'd19723: data <= 8'hFF;
            15'd19724: data <= 8'hFF;
            15'd19725: data <= 8'hFF;
            15'd19726: data <= 8'hFF;
            15'd19727: data <= 8'hFF;
            15'd19728: data <= 8'hFF;
            15'd19729: data <= 8'hFF;
            15'd19730: data <= 8'hFF;
            15'd19731: data <= 8'hFF;
            15'd19732: data <= 8'hFF;
            15'd19733: data <= 8'h03;
            15'd19734: data <= 8'h80;
            15'd19735: data <= 8'h00;
            15'd19736: data <= 8'h00;
            15'd19737: data <= 8'h00;
            15'd19738: data <= 8'h00;
            15'd19739: data <= 8'h00;
            15'd19740: data <= 8'h00;
            15'd19741: data <= 8'h00;
            15'd19742: data <= 8'h00;
            15'd19743: data <= 8'h00;
            15'd19744: data <= 8'h00;
            15'd19745: data <= 8'h03;
            15'd19746: data <= 8'hFF;
            15'd19747: data <= 8'hFF;
            15'd19748: data <= 8'hFF;
            15'd19749: data <= 8'hFC;
            15'd19750: data <= 8'h7F;
            15'd19751: data <= 8'hFF;
            15'd19752: data <= 8'h03;
            15'd19753: data <= 8'hFF;
            15'd19754: data <= 8'hFF;
            15'd19755: data <= 8'hFF;
            15'd19756: data <= 8'hFF;
            15'd19757: data <= 8'hFF;
            15'd19758: data <= 8'hFF;
            15'd19759: data <= 8'hFF;
            15'd19760: data <= 8'hFF;
            15'd19761: data <= 8'hFF;
            15'd19762: data <= 8'hFF;
            15'd19763: data <= 8'h01;
            15'd19764: data <= 8'h80;
            15'd19765: data <= 8'h00;
            15'd19766: data <= 8'h00;
            15'd19767: data <= 8'h00;
            15'd19768: data <= 8'h00;
            15'd19769: data <= 8'h00;
            15'd19770: data <= 8'h00;
            15'd19771: data <= 8'h00;
            15'd19772: data <= 8'h00;
            15'd19773: data <= 8'h00;
            15'd19774: data <= 8'h00;
            15'd19775: data <= 8'h03;
            15'd19776: data <= 8'hFF;
            15'd19777: data <= 8'hFF;
            15'd19778: data <= 8'hFF;
            15'd19779: data <= 8'hFC;
            15'd19780: data <= 8'h7F;
            15'd19781: data <= 8'hFF;
            15'd19782: data <= 8'h81;
            15'd19783: data <= 8'hFF;
            15'd19784: data <= 8'hFF;
            15'd19785: data <= 8'hFF;
            15'd19786: data <= 8'hFF;
            15'd19787: data <= 8'hFF;
            15'd19788: data <= 8'hFF;
            15'd19789: data <= 8'hFF;
            15'd19790: data <= 8'hFF;
            15'd19791: data <= 8'hFF;
            15'd19792: data <= 8'hFF;
            15'd19793: data <= 8'h81;
            15'd19794: data <= 8'h80;
            15'd19795: data <= 8'h00;
            15'd19796: data <= 8'h00;
            15'd19797: data <= 8'h00;
            15'd19798: data <= 8'h00;
            15'd19799: data <= 8'h00;
            15'd19800: data <= 8'h00;
            15'd19801: data <= 8'h00;
            15'd19802: data <= 8'h00;
            15'd19803: data <= 8'h00;
            15'd19804: data <= 8'h00;
            15'd19805: data <= 8'h03;
            15'd19806: data <= 8'hFF;
            15'd19807: data <= 8'hFF;
            15'd19808: data <= 8'hFF;
            15'd19809: data <= 8'hFC;
            15'd19810: data <= 8'h7F;
            15'd19811: data <= 8'hFF;
            15'd19812: data <= 8'hC1;
            15'd19813: data <= 8'hFF;
            15'd19814: data <= 8'hFF;
            15'd19815: data <= 8'hFF;
            15'd19816: data <= 8'hFF;
            15'd19817: data <= 8'hFF;
            15'd19818: data <= 8'hFF;
            15'd19819: data <= 8'hFF;
            15'd19820: data <= 8'hFF;
            15'd19821: data <= 8'hFF;
            15'd19822: data <= 8'hFF;
            15'd19823: data <= 8'h81;
            15'd19824: data <= 8'h80;
            15'd19825: data <= 8'h00;
            15'd19826: data <= 8'h00;
            15'd19827: data <= 8'h00;
            15'd19828: data <= 8'h00;
            15'd19829: data <= 8'h00;
            15'd19830: data <= 8'h00;
            15'd19831: data <= 8'h00;
            15'd19832: data <= 8'h00;
            15'd19833: data <= 8'h00;
            15'd19834: data <= 8'h00;
            15'd19835: data <= 8'h03;
            15'd19836: data <= 8'hFF;
            15'd19837: data <= 8'hFF;
            15'd19838: data <= 8'hFF;
            15'd19839: data <= 8'hF8;
            15'd19840: data <= 8'h7F;
            15'd19841: data <= 8'hFF;
            15'd19842: data <= 8'hE0;
            15'd19843: data <= 8'h7F;
            15'd19844: data <= 8'hFF;
            15'd19845: data <= 8'hFF;
            15'd19846: data <= 8'hFF;
            15'd19847: data <= 8'hFF;
            15'd19848: data <= 8'hFF;
            15'd19849: data <= 8'hFF;
            15'd19850: data <= 8'hFF;
            15'd19851: data <= 8'hFF;
            15'd19852: data <= 8'hFF;
            15'd19853: data <= 8'h81;
            15'd19854: data <= 8'h80;
            15'd19855: data <= 8'h00;
            15'd19856: data <= 8'h00;
            15'd19857: data <= 8'h00;
            15'd19858: data <= 8'h00;
            15'd19859: data <= 8'h00;
            15'd19860: data <= 8'h00;
            15'd19861: data <= 8'h00;
            15'd19862: data <= 8'h00;
            15'd19863: data <= 8'h00;
            15'd19864: data <= 8'h00;
            15'd19865: data <= 8'h03;
            15'd19866: data <= 8'hFF;
            15'd19867: data <= 8'hFF;
            15'd19868: data <= 8'hFF;
            15'd19869: data <= 8'hF0;
            15'd19870: data <= 8'h7F;
            15'd19871: data <= 8'hFF;
            15'd19872: data <= 8'hF0;
            15'd19873: data <= 8'h3F;
            15'd19874: data <= 8'hFF;
            15'd19875: data <= 8'hFF;
            15'd19876: data <= 8'hFF;
            15'd19877: data <= 8'hFF;
            15'd19878: data <= 8'hFF;
            15'd19879: data <= 8'hFF;
            15'd19880: data <= 8'hFF;
            15'd19881: data <= 8'hFF;
            15'd19882: data <= 8'hFF;
            15'd19883: data <= 8'h80;
            15'd19884: data <= 8'h80;
            15'd19885: data <= 8'h00;
            15'd19886: data <= 8'h00;
            15'd19887: data <= 8'h00;
            15'd19888: data <= 8'h00;
            15'd19889: data <= 8'h00;
            15'd19890: data <= 8'h00;
            15'd19891: data <= 8'h00;
            15'd19892: data <= 8'h00;
            15'd19893: data <= 8'h00;
            15'd19894: data <= 8'h00;
            15'd19895: data <= 8'h03;
            15'd19896: data <= 8'hFF;
            15'd19897: data <= 8'hFF;
            15'd19898: data <= 8'hFF;
            15'd19899: data <= 8'hF0;
            15'd19900: data <= 8'h7F;
            15'd19901: data <= 8'hFF;
            15'd19902: data <= 8'hF0;
            15'd19903: data <= 8'h1F;
            15'd19904: data <= 8'hFF;
            15'd19905: data <= 8'hFF;
            15'd19906: data <= 8'hFF;
            15'd19907: data <= 8'hFF;
            15'd19908: data <= 8'hFF;
            15'd19909: data <= 8'hFF;
            15'd19910: data <= 8'hFF;
            15'd19911: data <= 8'hFF;
            15'd19912: data <= 8'hFF;
            15'd19913: data <= 8'h80;
            15'd19914: data <= 8'h80;
            15'd19915: data <= 8'h00;
            15'd19916: data <= 8'h00;
            15'd19917: data <= 8'h00;
            15'd19918: data <= 8'h00;
            15'd19919: data <= 8'h00;
            15'd19920: data <= 8'h00;
            15'd19921: data <= 8'h00;
            15'd19922: data <= 8'h00;
            15'd19923: data <= 8'h00;
            15'd19924: data <= 8'h00;
            15'd19925: data <= 8'h03;
            15'd19926: data <= 8'hFF;
            15'd19927: data <= 8'hFF;
            15'd19928: data <= 8'hFF;
            15'd19929: data <= 8'hF0;
            15'd19930: data <= 8'h3F;
            15'd19931: data <= 8'hFF;
            15'd19932: data <= 8'hF8;
            15'd19933: data <= 8'h07;
            15'd19934: data <= 8'hFF;
            15'd19935: data <= 8'hFF;
            15'd19936: data <= 8'hFF;
            15'd19937: data <= 8'hFF;
            15'd19938: data <= 8'hFF;
            15'd19939: data <= 8'hFF;
            15'd19940: data <= 8'hFF;
            15'd19941: data <= 8'hFF;
            15'd19942: data <= 8'hFF;
            15'd19943: data <= 8'h80;
            15'd19944: data <= 8'h80;
            15'd19945: data <= 8'h00;
            15'd19946: data <= 8'h00;
            15'd19947: data <= 8'h00;
            15'd19948: data <= 8'h00;
            15'd19949: data <= 8'h00;
            15'd19950: data <= 8'h00;
            15'd19951: data <= 8'h00;
            15'd19952: data <= 8'h00;
            15'd19953: data <= 8'h00;
            15'd19954: data <= 8'h00;
            15'd19955: data <= 8'h03;
            15'd19956: data <= 8'hFF;
            15'd19957: data <= 8'hFF;
            15'd19958: data <= 8'hFF;
            15'd19959: data <= 8'hF8;
            15'd19960: data <= 8'h3F;
            15'd19961: data <= 8'hFF;
            15'd19962: data <= 8'hFE;
            15'd19963: data <= 8'h01;
            15'd19964: data <= 8'hFF;
            15'd19965: data <= 8'hFF;
            15'd19966: data <= 8'hFF;
            15'd19967: data <= 8'hFF;
            15'd19968: data <= 8'hFF;
            15'd19969: data <= 8'hFF;
            15'd19970: data <= 8'hFF;
            15'd19971: data <= 8'hFF;
            15'd19972: data <= 8'hFF;
            15'd19973: data <= 8'hC0;
            15'd19974: data <= 8'h00;
            15'd19975: data <= 8'h00;
            15'd19976: data <= 8'h00;
            15'd19977: data <= 8'h00;
            15'd19978: data <= 8'h00;
            15'd19979: data <= 8'h00;
            15'd19980: data <= 8'h00;
            15'd19981: data <= 8'h00;
            15'd19982: data <= 8'h00;
            15'd19983: data <= 8'h00;
            15'd19984: data <= 8'h00;
            15'd19985: data <= 8'h03;
            15'd19986: data <= 8'hFF;
            15'd19987: data <= 8'hFF;
            15'd19988: data <= 8'hFF;
            15'd19989: data <= 8'hF8;
            15'd19990: data <= 8'h3F;
            15'd19991: data <= 8'hFF;
            15'd19992: data <= 8'hFF;
            15'd19993: data <= 8'h00;
            15'd19994: data <= 8'hFF;
            15'd19995: data <= 8'hFF;
            15'd19996: data <= 8'hFF;
            15'd19997: data <= 8'hFF;
            15'd19998: data <= 8'hFF;
            15'd19999: data <= 8'hFF;
            15'd20000: data <= 8'hFF;
            15'd20001: data <= 8'hFF;
            15'd20002: data <= 8'hFF;
            15'd20003: data <= 8'hC0;
            15'd20004: data <= 8'h00;
            15'd20005: data <= 8'h00;
            15'd20006: data <= 8'h00;
            15'd20007: data <= 8'h00;
            15'd20008: data <= 8'h00;
            15'd20009: data <= 8'h00;
            15'd20010: data <= 8'h00;
            15'd20011: data <= 8'h00;
            15'd20012: data <= 8'h00;
            15'd20013: data <= 8'h00;
            15'd20014: data <= 8'h00;
            15'd20015: data <= 8'h03;
            15'd20016: data <= 8'hFF;
            15'd20017: data <= 8'hFF;
            15'd20018: data <= 8'hFF;
            15'd20019: data <= 8'hF8;
            15'd20020: data <= 8'h7F;
            15'd20021: data <= 8'hFF;
            15'd20022: data <= 8'hFF;
            15'd20023: data <= 8'h80;
            15'd20024: data <= 8'h1F;
            15'd20025: data <= 8'hFF;
            15'd20026: data <= 8'hFF;
            15'd20027: data <= 8'hFF;
            15'd20028: data <= 8'hFF;
            15'd20029: data <= 8'hFF;
            15'd20030: data <= 8'hFF;
            15'd20031: data <= 8'hFF;
            15'd20032: data <= 8'hFF;
            15'd20033: data <= 8'hC0;
            15'd20034: data <= 8'h00;
            15'd20035: data <= 8'h00;
            15'd20036: data <= 8'h00;
            15'd20037: data <= 8'h00;
            15'd20038: data <= 8'h00;
            15'd20039: data <= 8'h00;
            15'd20040: data <= 8'h00;
            15'd20041: data <= 8'h00;
            15'd20042: data <= 8'h00;
            15'd20043: data <= 8'h00;
            15'd20044: data <= 8'h00;
            15'd20045: data <= 8'h03;
            15'd20046: data <= 8'hFF;
            15'd20047: data <= 8'hFF;
            15'd20048: data <= 8'hFF;
            15'd20049: data <= 8'hF8;
            15'd20050: data <= 8'h7F;
            15'd20051: data <= 8'hFF;
            15'd20052: data <= 8'hFF;
            15'd20053: data <= 8'hC0;
            15'd20054: data <= 8'h07;
            15'd20055: data <= 8'hFF;
            15'd20056: data <= 8'hFF;
            15'd20057: data <= 8'hFF;
            15'd20058: data <= 8'hFF;
            15'd20059: data <= 8'hFF;
            15'd20060: data <= 8'hFF;
            15'd20061: data <= 8'hFF;
            15'd20062: data <= 8'hFF;
            15'd20063: data <= 8'hC0;
            15'd20064: data <= 8'h00;
            15'd20065: data <= 8'h00;
            15'd20066: data <= 8'h00;
            15'd20067: data <= 8'h00;
            15'd20068: data <= 8'h00;
            15'd20069: data <= 8'h00;
            15'd20070: data <= 8'h00;
            15'd20071: data <= 8'h00;
            15'd20072: data <= 8'h00;
            15'd20073: data <= 8'h00;
            15'd20074: data <= 8'h00;
            15'd20075: data <= 8'h03;
            15'd20076: data <= 8'hFF;
            15'd20077: data <= 8'hFF;
            15'd20078: data <= 8'hFF;
            15'd20079: data <= 8'hF8;
            15'd20080: data <= 8'h7F;
            15'd20081: data <= 8'hFF;
            15'd20082: data <= 8'hFF;
            15'd20083: data <= 8'hE0;
            15'd20084: data <= 8'h01;
            15'd20085: data <= 8'hFF;
            15'd20086: data <= 8'hFF;
            15'd20087: data <= 8'hFF;
            15'd20088: data <= 8'hFF;
            15'd20089: data <= 8'hFF;
            15'd20090: data <= 8'hFF;
            15'd20091: data <= 8'hFF;
            15'd20092: data <= 8'hFF;
            15'd20093: data <= 8'hC0;
            15'd20094: data <= 8'h00;
            15'd20095: data <= 8'h00;
            15'd20096: data <= 8'h00;
            15'd20097: data <= 8'h00;
            15'd20098: data <= 8'h00;
            15'd20099: data <= 8'h00;
            15'd20100: data <= 8'h00;
            15'd20101: data <= 8'h00;
            15'd20102: data <= 8'h00;
            15'd20103: data <= 8'h00;
            15'd20104: data <= 8'h00;
            15'd20105: data <= 8'h03;
            15'd20106: data <= 8'hFF;
            15'd20107: data <= 8'hFF;
            15'd20108: data <= 8'hFF;
            15'd20109: data <= 8'hF8;
            15'd20110: data <= 8'h7F;
            15'd20111: data <= 8'hFF;
            15'd20112: data <= 8'hFF;
            15'd20113: data <= 8'hF8;
            15'd20114: data <= 8'h00;
            15'd20115: data <= 8'h7F;
            15'd20116: data <= 8'hFC;
            15'd20117: data <= 8'h7F;
            15'd20118: data <= 8'hFF;
            15'd20119: data <= 8'hFF;
            15'd20120: data <= 8'hFF;
            15'd20121: data <= 8'hFF;
            15'd20122: data <= 8'hFF;
            15'd20123: data <= 8'hE0;
            15'd20124: data <= 8'h00;
            15'd20125: data <= 8'h00;
            15'd20126: data <= 8'h00;
            15'd20127: data <= 8'h00;
            15'd20128: data <= 8'h00;
            15'd20129: data <= 8'h00;
            15'd20130: data <= 8'h00;
            15'd20131: data <= 8'h00;
            15'd20132: data <= 8'h00;
            15'd20133: data <= 8'h00;
            15'd20134: data <= 8'h00;
            15'd20135: data <= 8'h03;
            15'd20136: data <= 8'hFF;
            15'd20137: data <= 8'hFF;
            15'd20138: data <= 8'hFF;
            15'd20139: data <= 8'hF8;
            15'd20140: data <= 8'h7F;
            15'd20141: data <= 8'hFF;
            15'd20142: data <= 8'hFF;
            15'd20143: data <= 8'hFC;
            15'd20144: data <= 8'h00;
            15'd20145: data <= 8'h00;
            15'd20146: data <= 8'hC0;
            15'd20147: data <= 8'h3F;
            15'd20148: data <= 8'hFF;
            15'd20149: data <= 8'hFF;
            15'd20150: data <= 8'hFF;
            15'd20151: data <= 8'hFF;
            15'd20152: data <= 8'hFF;
            15'd20153: data <= 8'hE0;
            15'd20154: data <= 8'h00;
            15'd20155: data <= 8'h00;
            15'd20156: data <= 8'h00;
            15'd20157: data <= 8'h00;
            15'd20158: data <= 8'h00;
            15'd20159: data <= 8'h00;
            15'd20160: data <= 8'h00;
            15'd20161: data <= 8'h00;
            15'd20162: data <= 8'h00;
            15'd20163: data <= 8'h00;
            15'd20164: data <= 8'h00;
            15'd20165: data <= 8'h03;
            15'd20166: data <= 8'hFF;
            15'd20167: data <= 8'hFF;
            15'd20168: data <= 8'hFF;
            15'd20169: data <= 8'hF0;
            15'd20170: data <= 8'h7F;
            15'd20171: data <= 8'hFF;
            15'd20172: data <= 8'hFF;
            15'd20173: data <= 8'hFF;
            15'd20174: data <= 8'h00;
            15'd20175: data <= 8'h00;
            15'd20176: data <= 8'h00;
            15'd20177: data <= 8'h1F;
            15'd20178: data <= 8'hFF;
            15'd20179: data <= 8'hFF;
            15'd20180: data <= 8'hFF;
            15'd20181: data <= 8'hFF;
            15'd20182: data <= 8'hFF;
            15'd20183: data <= 8'hE0;
            15'd20184: data <= 8'h00;
            15'd20185: data <= 8'h00;
            15'd20186: data <= 8'h00;
            15'd20187: data <= 8'h00;
            15'd20188: data <= 8'h00;
            15'd20189: data <= 8'h00;
            15'd20190: data <= 8'h00;
            15'd20191: data <= 8'h00;
            15'd20192: data <= 8'h00;
            15'd20193: data <= 8'h00;
            15'd20194: data <= 8'h00;
            15'd20195: data <= 8'h03;
            15'd20196: data <= 8'hFF;
            15'd20197: data <= 8'hFF;
            15'd20198: data <= 8'hFF;
            15'd20199: data <= 8'hF0;
            15'd20200: data <= 8'h7F;
            15'd20201: data <= 8'hFF;
            15'd20202: data <= 8'hFF;
            15'd20203: data <= 8'hFF;
            15'd20204: data <= 8'hC0;
            15'd20205: data <= 8'h00;
            15'd20206: data <= 8'h00;
            15'd20207: data <= 8'h3F;
            15'd20208: data <= 8'hFF;
            15'd20209: data <= 8'hFF;
            15'd20210: data <= 8'hFF;
            15'd20211: data <= 8'hFF;
            15'd20212: data <= 8'hFF;
            15'd20213: data <= 8'hE0;
            15'd20214: data <= 8'h00;
            15'd20215: data <= 8'h00;
            15'd20216: data <= 8'h00;
            15'd20217: data <= 8'h00;
            15'd20218: data <= 8'h00;
            15'd20219: data <= 8'h00;
            15'd20220: data <= 8'h00;
            15'd20221: data <= 8'h00;
            15'd20222: data <= 8'h00;
            15'd20223: data <= 8'h00;
            15'd20224: data <= 8'h00;
            15'd20225: data <= 8'h03;
            15'd20226: data <= 8'hFF;
            15'd20227: data <= 8'hFF;
            15'd20228: data <= 8'hFF;
            15'd20229: data <= 8'hF0;
            15'd20230: data <= 8'h7F;
            15'd20231: data <= 8'hFF;
            15'd20232: data <= 8'hFF;
            15'd20233: data <= 8'hFF;
            15'd20234: data <= 8'hF0;
            15'd20235: data <= 8'h00;
            15'd20236: data <= 8'h00;
            15'd20237: data <= 8'h3F;
            15'd20238: data <= 8'hFF;
            15'd20239: data <= 8'hFF;
            15'd20240: data <= 8'hFF;
            15'd20241: data <= 8'hFF;
            15'd20242: data <= 8'hFF;
            15'd20243: data <= 8'hE0;
            15'd20244: data <= 8'h00;
            15'd20245: data <= 8'h00;
            15'd20246: data <= 8'h00;
            15'd20247: data <= 8'h00;
            15'd20248: data <= 8'h00;
            15'd20249: data <= 8'h00;
            15'd20250: data <= 8'h00;
            15'd20251: data <= 8'h00;
            15'd20252: data <= 8'h00;
            15'd20253: data <= 8'h00;
            15'd20254: data <= 8'h00;
            15'd20255: data <= 8'h03;
            15'd20256: data <= 8'hFF;
            15'd20257: data <= 8'hFF;
            15'd20258: data <= 8'hFF;
            15'd20259: data <= 8'hF0;
            15'd20260: data <= 8'h7F;
            15'd20261: data <= 8'hFF;
            15'd20262: data <= 8'hFF;
            15'd20263: data <= 8'hFF;
            15'd20264: data <= 8'hF8;
            15'd20265: data <= 8'h00;
            15'd20266: data <= 8'h00;
            15'd20267: data <= 8'h7F;
            15'd20268: data <= 8'hFF;
            15'd20269: data <= 8'hFF;
            15'd20270: data <= 8'hFF;
            15'd20271: data <= 8'hFF;
            15'd20272: data <= 8'hFF;
            15'd20273: data <= 8'hE0;
            15'd20274: data <= 8'h00;
            15'd20275: data <= 8'h00;
            15'd20276: data <= 8'h00;
            15'd20277: data <= 8'h00;
            15'd20278: data <= 8'h00;
            15'd20279: data <= 8'h00;
            15'd20280: data <= 8'h00;
            15'd20281: data <= 8'h00;
            15'd20282: data <= 8'h00;
            15'd20283: data <= 8'h00;
            15'd20284: data <= 8'h00;
            15'd20285: data <= 8'h03;
            15'd20286: data <= 8'hFF;
            15'd20287: data <= 8'hFF;
            15'd20288: data <= 8'hFF;
            15'd20289: data <= 8'hF0;
            15'd20290: data <= 8'h7F;
            15'd20291: data <= 8'hFF;
            15'd20292: data <= 8'hFF;
            15'd20293: data <= 8'hFF;
            15'd20294: data <= 8'hFF;
            15'd20295: data <= 8'hC0;
            15'd20296: data <= 8'h03;
            15'd20297: data <= 8'hFF;
            15'd20298: data <= 8'hFF;
            15'd20299: data <= 8'hFF;
            15'd20300: data <= 8'hFF;
            15'd20301: data <= 8'hFF;
            15'd20302: data <= 8'hFF;
            15'd20303: data <= 8'hF0;
            15'd20304: data <= 8'h00;
            15'd20305: data <= 8'h00;
            15'd20306: data <= 8'h00;
            15'd20307: data <= 8'h00;
            15'd20308: data <= 8'h00;
            15'd20309: data <= 8'h00;
            15'd20310: data <= 8'h00;
            15'd20311: data <= 8'h00;
            15'd20312: data <= 8'h00;
            15'd20313: data <= 8'h00;
            15'd20314: data <= 8'h00;
            15'd20315: data <= 8'h03;
            15'd20316: data <= 8'hFF;
            15'd20317: data <= 8'hFF;
            15'd20318: data <= 8'hFF;
            15'd20319: data <= 8'hF0;
            15'd20320: data <= 8'h7F;
            15'd20321: data <= 8'hFF;
            15'd20322: data <= 8'hFF;
            15'd20323: data <= 8'hFF;
            15'd20324: data <= 8'hFF;
            15'd20325: data <= 8'hFF;
            15'd20326: data <= 8'hFF;
            15'd20327: data <= 8'hFF;
            15'd20328: data <= 8'hFF;
            15'd20329: data <= 8'hFF;
            15'd20330: data <= 8'hFF;
            15'd20331: data <= 8'hFF;
            15'd20332: data <= 8'hFF;
            15'd20333: data <= 8'hF0;
            15'd20334: data <= 8'h00;
            15'd20335: data <= 8'h00;
            15'd20336: data <= 8'h00;
            15'd20337: data <= 8'h00;
            15'd20338: data <= 8'h00;
            15'd20339: data <= 8'h00;
            15'd20340: data <= 8'h00;
            15'd20341: data <= 8'h00;
            15'd20342: data <= 8'h00;
            15'd20343: data <= 8'h00;
            15'd20344: data <= 8'h00;
            15'd20345: data <= 8'h03;
            15'd20346: data <= 8'hFF;
            15'd20347: data <= 8'hFF;
            15'd20348: data <= 8'hFF;
            15'd20349: data <= 8'hF0;
            15'd20350: data <= 8'h7F;
            15'd20351: data <= 8'hFF;
            15'd20352: data <= 8'hFF;
            15'd20353: data <= 8'hFF;
            15'd20354: data <= 8'hFF;
            15'd20355: data <= 8'hFF;
            15'd20356: data <= 8'hFF;
            15'd20357: data <= 8'hFF;
            15'd20358: data <= 8'hFF;
            15'd20359: data <= 8'hFF;
            15'd20360: data <= 8'hFF;
            15'd20361: data <= 8'hFF;
            15'd20362: data <= 8'hFF;
            15'd20363: data <= 8'hF0;
            15'd20364: data <= 8'h00;
            15'd20365: data <= 8'h00;
            15'd20366: data <= 8'h00;
            15'd20367: data <= 8'h00;
            15'd20368: data <= 8'h00;
            15'd20369: data <= 8'h00;
            15'd20370: data <= 8'h00;
            15'd20371: data <= 8'h00;
            15'd20372: data <= 8'h00;
            15'd20373: data <= 8'h00;
            15'd20374: data <= 8'h00;
            15'd20375: data <= 8'h03;
            15'd20376: data <= 8'hFF;
            15'd20377: data <= 8'hFF;
            15'd20378: data <= 8'hFF;
            15'd20379: data <= 8'hF0;
            15'd20380: data <= 8'h7F;
            15'd20381: data <= 8'hFF;
            15'd20382: data <= 8'hFF;
            15'd20383: data <= 8'hFF;
            15'd20384: data <= 8'hFF;
            15'd20385: data <= 8'hFF;
            15'd20386: data <= 8'hFF;
            15'd20387: data <= 8'hFF;
            15'd20388: data <= 8'hFF;
            15'd20389: data <= 8'hFF;
            15'd20390: data <= 8'hFF;
            15'd20391: data <= 8'hFF;
            15'd20392: data <= 8'hFF;
            15'd20393: data <= 8'hF0;
            15'd20394: data <= 8'h00;
            15'd20395: data <= 8'h00;
            15'd20396: data <= 8'h00;
            15'd20397: data <= 8'h00;
            15'd20398: data <= 8'h00;
            15'd20399: data <= 8'h00;
            15'd20400: data <= 8'h00;
            15'd20401: data <= 8'h00;
            15'd20402: data <= 8'h00;
            15'd20403: data <= 8'h00;
            15'd20404: data <= 8'h00;
            15'd20405: data <= 8'h03;
            15'd20406: data <= 8'hFF;
            15'd20407: data <= 8'hFF;
            15'd20408: data <= 8'hFF;
            15'd20409: data <= 8'hF0;
            15'd20410: data <= 8'h7F;
            15'd20411: data <= 8'hFF;
            15'd20412: data <= 8'hFF;
            15'd20413: data <= 8'hFF;
            15'd20414: data <= 8'hFF;
            15'd20415: data <= 8'hFF;
            15'd20416: data <= 8'hFF;
            15'd20417: data <= 8'hFF;
            15'd20418: data <= 8'hFF;
            15'd20419: data <= 8'hFF;
            15'd20420: data <= 8'hFF;
            15'd20421: data <= 8'hFF;
            15'd20422: data <= 8'hFF;
            15'd20423: data <= 8'hF0;
            15'd20424: data <= 8'h00;
            15'd20425: data <= 8'h00;
            15'd20426: data <= 8'h00;
            15'd20427: data <= 8'h00;
            15'd20428: data <= 8'h00;
            15'd20429: data <= 8'h00;
            15'd20430: data <= 8'h00;
            15'd20431: data <= 8'h00;
            15'd20432: data <= 8'h00;
            15'd20433: data <= 8'h00;
            15'd20434: data <= 8'h00;
            15'd20435: data <= 8'h03;
            15'd20436: data <= 8'hFF;
            15'd20437: data <= 8'hFF;
            15'd20438: data <= 8'hFF;
            15'd20439: data <= 8'hF0;
            15'd20440: data <= 8'h7F;
            15'd20441: data <= 8'hFF;
            15'd20442: data <= 8'hFF;
            15'd20443: data <= 8'hFF;
            15'd20444: data <= 8'hFF;
            15'd20445: data <= 8'hFF;
            15'd20446: data <= 8'hFF;
            15'd20447: data <= 8'hFF;
            15'd20448: data <= 8'hFF;
            15'd20449: data <= 8'hFF;
            15'd20450: data <= 8'hFF;
            15'd20451: data <= 8'hFF;
            15'd20452: data <= 8'hFF;
            15'd20453: data <= 8'hF0;
            15'd20454: data <= 8'h00;
            15'd20455: data <= 8'h00;
            15'd20456: data <= 8'h00;
            15'd20457: data <= 8'h00;
            15'd20458: data <= 8'h00;
            15'd20459: data <= 8'h00;
            15'd20460: data <= 8'h00;
            15'd20461: data <= 8'h00;
            15'd20462: data <= 8'h00;
            15'd20463: data <= 8'h00;
            15'd20464: data <= 8'h00;
            15'd20465: data <= 8'h03;
            15'd20466: data <= 8'hFF;
            15'd20467: data <= 8'hFF;
            15'd20468: data <= 8'hFF;
            15'd20469: data <= 8'hF0;
            15'd20470: data <= 8'h7F;
            15'd20471: data <= 8'hFF;
            15'd20472: data <= 8'hFF;
            15'd20473: data <= 8'hFF;
            15'd20474: data <= 8'hFF;
            15'd20475: data <= 8'hFF;
            15'd20476: data <= 8'hFF;
            15'd20477: data <= 8'hFF;
            15'd20478: data <= 8'hFF;
            15'd20479: data <= 8'hFF;
            15'd20480: data <= 8'hFF;
            15'd20481: data <= 8'hFF;
            15'd20482: data <= 8'hFF;
            15'd20483: data <= 8'hF8;
            15'd20484: data <= 8'h00;
            15'd20485: data <= 8'h00;
            15'd20486: data <= 8'h00;
            15'd20487: data <= 8'h00;
            15'd20488: data <= 8'h00;
            15'd20489: data <= 8'h00;
            15'd20490: data <= 8'h00;
            15'd20491: data <= 8'h00;
            15'd20492: data <= 8'h00;
            15'd20493: data <= 8'h00;
            15'd20494: data <= 8'h00;
            15'd20495: data <= 8'h03;
            15'd20496: data <= 8'hFF;
            15'd20497: data <= 8'hFF;
            15'd20498: data <= 8'hFF;
            15'd20499: data <= 8'hE0;
            15'd20500: data <= 8'h7F;
            15'd20501: data <= 8'hFF;
            15'd20502: data <= 8'hFF;
            15'd20503: data <= 8'hFF;
            15'd20504: data <= 8'hFF;
            15'd20505: data <= 8'hFF;
            15'd20506: data <= 8'hFF;
            15'd20507: data <= 8'hFF;
            15'd20508: data <= 8'hFF;
            15'd20509: data <= 8'hFF;
            15'd20510: data <= 8'hFF;
            15'd20511: data <= 8'hFF;
            15'd20512: data <= 8'hFF;
            15'd20513: data <= 8'hF8;
            15'd20514: data <= 8'h00;
            15'd20515: data <= 8'h00;
            15'd20516: data <= 8'h00;
            15'd20517: data <= 8'h00;
            15'd20518: data <= 8'h00;
            15'd20519: data <= 8'h00;
            15'd20520: data <= 8'h00;
            15'd20521: data <= 8'h00;
            15'd20522: data <= 8'h00;
            15'd20523: data <= 8'h00;
            15'd20524: data <= 8'h00;
            15'd20525: data <= 8'h03;
            15'd20526: data <= 8'hFF;
            15'd20527: data <= 8'hFF;
            15'd20528: data <= 8'hFF;
            15'd20529: data <= 8'hE0;
            15'd20530: data <= 8'h7F;
            15'd20531: data <= 8'hFF;
            15'd20532: data <= 8'hFF;
            15'd20533: data <= 8'hFF;
            15'd20534: data <= 8'hFF;
            15'd20535: data <= 8'hFF;
            15'd20536: data <= 8'hFF;
            15'd20537: data <= 8'hFF;
            15'd20538: data <= 8'hFF;
            15'd20539: data <= 8'hFF;
            15'd20540: data <= 8'hFF;
            15'd20541: data <= 8'hFF;
            15'd20542: data <= 8'hFF;
            15'd20543: data <= 8'hF8;
            15'd20544: data <= 8'h00;
            15'd20545: data <= 8'h00;
            15'd20546: data <= 8'h00;
            15'd20547: data <= 8'h00;
            15'd20548: data <= 8'h00;
            15'd20549: data <= 8'h00;
            15'd20550: data <= 8'h00;
            15'd20551: data <= 8'h00;
            15'd20552: data <= 8'h00;
            15'd20553: data <= 8'h00;
            15'd20554: data <= 8'h00;
            15'd20555: data <= 8'h03;
            15'd20556: data <= 8'hFF;
            15'd20557: data <= 8'hFF;
            15'd20558: data <= 8'hFF;
            15'd20559: data <= 8'hE0;
            15'd20560: data <= 8'h7F;
            15'd20561: data <= 8'hFF;
            15'd20562: data <= 8'hFF;
            15'd20563: data <= 8'hFF;
            15'd20564: data <= 8'hFF;
            15'd20565: data <= 8'hFF;
            15'd20566: data <= 8'hFF;
            15'd20567: data <= 8'hFF;
            15'd20568: data <= 8'hFF;
            15'd20569: data <= 8'hFF;
            15'd20570: data <= 8'hFF;
            15'd20571: data <= 8'hFF;
            15'd20572: data <= 8'hFF;
            15'd20573: data <= 8'hF8;
            15'd20574: data <= 8'h00;
            15'd20575: data <= 8'h00;
            15'd20576: data <= 8'h00;
            15'd20577: data <= 8'h00;
            15'd20578: data <= 8'h00;
            15'd20579: data <= 8'h00;
            15'd20580: data <= 8'h00;
            15'd20581: data <= 8'h00;
            15'd20582: data <= 8'h00;
            15'd20583: data <= 8'h00;
            15'd20584: data <= 8'h00;
            15'd20585: data <= 8'h03;
            15'd20586: data <= 8'hFF;
            15'd20587: data <= 8'hFF;
            15'd20588: data <= 8'hFF;
            15'd20589: data <= 8'hE0;
            15'd20590: data <= 8'h7F;
            15'd20591: data <= 8'hFF;
            15'd20592: data <= 8'hFF;
            15'd20593: data <= 8'hFF;
            15'd20594: data <= 8'hFF;
            15'd20595: data <= 8'hFF;
            15'd20596: data <= 8'hFF;
            15'd20597: data <= 8'hFF;
            15'd20598: data <= 8'hFF;
            15'd20599: data <= 8'hFF;
            15'd20600: data <= 8'hFF;
            15'd20601: data <= 8'hFF;
            15'd20602: data <= 8'hFF;
            15'd20603: data <= 8'hF8;
            15'd20604: data <= 8'h00;
            15'd20605: data <= 8'h00;
            15'd20606: data <= 8'h00;
            15'd20607: data <= 8'h00;
            15'd20608: data <= 8'h00;
            15'd20609: data <= 8'h00;
            15'd20610: data <= 8'h00;
            15'd20611: data <= 8'h00;
            15'd20612: data <= 8'h00;
            15'd20613: data <= 8'h00;
            15'd20614: data <= 8'h00;
            15'd20615: data <= 8'h03;
            15'd20616: data <= 8'hFF;
            15'd20617: data <= 8'hFF;
            15'd20618: data <= 8'hFF;
            15'd20619: data <= 8'hF0;
            15'd20620: data <= 8'hFF;
            15'd20621: data <= 8'hFF;
            15'd20622: data <= 8'hFF;
            15'd20623: data <= 8'hFF;
            15'd20624: data <= 8'hFF;
            15'd20625: data <= 8'hFF;
            15'd20626: data <= 8'hFF;
            15'd20627: data <= 8'hFF;
            15'd20628: data <= 8'hFF;
            15'd20629: data <= 8'hFF;
            15'd20630: data <= 8'hFF;
            15'd20631: data <= 8'hFF;
            15'd20632: data <= 8'hFF;
            15'd20633: data <= 8'hFC;
            15'd20634: data <= 8'h00;
            15'd20635: data <= 8'h00;
            15'd20636: data <= 8'h00;
            15'd20637: data <= 8'h00;
            15'd20638: data <= 8'h00;
            15'd20639: data <= 8'h00;
            15'd20640: data <= 8'h00;
            15'd20641: data <= 8'h00;
            15'd20642: data <= 8'h00;
            15'd20643: data <= 8'h00;
            15'd20644: data <= 8'h00;
            15'd20645: data <= 8'h03;
            15'd20646: data <= 8'hFF;
            15'd20647: data <= 8'hFF;
            15'd20648: data <= 8'hFF;
            15'd20649: data <= 8'hFF;
            15'd20650: data <= 8'hFF;
            15'd20651: data <= 8'hFF;
            15'd20652: data <= 8'hFF;
            15'd20653: data <= 8'hFF;
            15'd20654: data <= 8'hFF;
            15'd20655: data <= 8'hFF;
            15'd20656: data <= 8'hFF;
            15'd20657: data <= 8'hFF;
            15'd20658: data <= 8'hFF;
            15'd20659: data <= 8'hFF;
            15'd20660: data <= 8'hFF;
            15'd20661: data <= 8'hFF;
            15'd20662: data <= 8'hFF;
            15'd20663: data <= 8'hFF;
            15'd20664: data <= 8'h80;
            15'd20665: data <= 8'h00;
            15'd20666: data <= 8'h00;
            15'd20667: data <= 8'h00;
            15'd20668: data <= 8'h00;
            15'd20669: data <= 8'h00;
            15'd20670: data <= 8'h00;
            15'd20671: data <= 8'h00;
            15'd20672: data <= 8'h00;
            15'd20673: data <= 8'h00;
            15'd20674: data <= 8'h00;
            15'd20675: data <= 8'h03;
            15'd20676: data <= 8'hFF;
            15'd20677: data <= 8'hFF;
            15'd20678: data <= 8'hFF;
            15'd20679: data <= 8'hFF;
            15'd20680: data <= 8'hFF;
            15'd20681: data <= 8'hFF;
            15'd20682: data <= 8'hFF;
            15'd20683: data <= 8'hFF;
            15'd20684: data <= 8'hFF;
            15'd20685: data <= 8'hFF;
            15'd20686: data <= 8'hFF;
            15'd20687: data <= 8'hFF;
            15'd20688: data <= 8'hFF;
            15'd20689: data <= 8'hFF;
            15'd20690: data <= 8'hFF;
            15'd20691: data <= 8'hFF;
            15'd20692: data <= 8'hFF;
            15'd20693: data <= 8'hFF;
            15'd20694: data <= 8'h80;
            15'd20695: data <= 8'h00;
            15'd20696: data <= 8'h00;
            15'd20697: data <= 8'h00;
            15'd20698: data <= 8'h00;
            15'd20699: data <= 8'h00;
            15'd20700: data <= 8'h00;
            15'd20701: data <= 8'h00;
            15'd20702: data <= 8'h00;
            15'd20703: data <= 8'h00;
            15'd20704: data <= 8'h00;
            15'd20705: data <= 8'h03;
            15'd20706: data <= 8'hFF;
            15'd20707: data <= 8'hFF;
            15'd20708: data <= 8'hFF;
            15'd20709: data <= 8'hFF;
            15'd20710: data <= 8'hFF;
            15'd20711: data <= 8'hFF;
            15'd20712: data <= 8'hFF;
            15'd20713: data <= 8'hFF;
            15'd20714: data <= 8'hFF;
            15'd20715: data <= 8'hFF;
            15'd20716: data <= 8'hFF;
            15'd20717: data <= 8'hFF;
            15'd20718: data <= 8'hFF;
            15'd20719: data <= 8'hFF;
            15'd20720: data <= 8'hFF;
            15'd20721: data <= 8'hFF;
            15'd20722: data <= 8'hFF;
            15'd20723: data <= 8'hFF;
            15'd20724: data <= 8'h80;
            15'd20725: data <= 8'h00;
            15'd20726: data <= 8'h00;
            15'd20727: data <= 8'h00;
            15'd20728: data <= 8'h00;
            15'd20729: data <= 8'h00;
            15'd20730: data <= 8'h00;
            15'd20731: data <= 8'h00;
            15'd20732: data <= 8'h00;
            15'd20733: data <= 8'h00;
            15'd20734: data <= 8'h00;
            15'd20735: data <= 8'h03;
            15'd20736: data <= 8'hFF;
            15'd20737: data <= 8'hFF;
            15'd20738: data <= 8'hFF;
            15'd20739: data <= 8'hFF;
            15'd20740: data <= 8'hFF;
            15'd20741: data <= 8'hFF;
            15'd20742: data <= 8'hFF;
            15'd20743: data <= 8'hFF;
            15'd20744: data <= 8'hFF;
            15'd20745: data <= 8'hFF;
            15'd20746: data <= 8'hFF;
            15'd20747: data <= 8'hFF;
            15'd20748: data <= 8'hFF;
            15'd20749: data <= 8'hFF;
            15'd20750: data <= 8'hFF;
            15'd20751: data <= 8'hFF;
            15'd20752: data <= 8'hFF;
            15'd20753: data <= 8'hFF;
            15'd20754: data <= 8'h80;
            15'd20755: data <= 8'h00;
            15'd20756: data <= 8'h00;
            15'd20757: data <= 8'h00;
            15'd20758: data <= 8'h00;
            15'd20759: data <= 8'h00;
            15'd20760: data <= 8'h00;
            15'd20761: data <= 8'h00;
            15'd20762: data <= 8'h00;
            15'd20763: data <= 8'h00;
            15'd20764: data <= 8'h00;
            15'd20765: data <= 8'h03;
            15'd20766: data <= 8'hFF;
            15'd20767: data <= 8'hFF;
            15'd20768: data <= 8'hFF;
            15'd20769: data <= 8'hFF;
            15'd20770: data <= 8'hFF;
            15'd20771: data <= 8'hFF;
            15'd20772: data <= 8'hFF;
            15'd20773: data <= 8'hFF;
            15'd20774: data <= 8'hFF;
            15'd20775: data <= 8'hFF;
            15'd20776: data <= 8'hFF;
            15'd20777: data <= 8'hFF;
            15'd20778: data <= 8'hFF;
            15'd20779: data <= 8'hFF;
            15'd20780: data <= 8'hFF;
            15'd20781: data <= 8'hFF;
            15'd20782: data <= 8'hFF;
            15'd20783: data <= 8'hFF;
            15'd20784: data <= 8'h80;
            15'd20785: data <= 8'h00;
            15'd20786: data <= 8'h00;
            15'd20787: data <= 8'h00;
            15'd20788: data <= 8'h00;
            15'd20789: data <= 8'h00;
            15'd20790: data <= 8'h00;
            15'd20791: data <= 8'h00;
            15'd20792: data <= 8'h00;
            15'd20793: data <= 8'h00;
            15'd20794: data <= 8'h00;
            15'd20795: data <= 8'h03;
            15'd20796: data <= 8'hFF;
            15'd20797: data <= 8'hFF;
            15'd20798: data <= 8'hFF;
            15'd20799: data <= 8'hFF;
            15'd20800: data <= 8'hFF;
            15'd20801: data <= 8'hFF;
            15'd20802: data <= 8'hFF;
            15'd20803: data <= 8'hFF;
            15'd20804: data <= 8'hFF;
            15'd20805: data <= 8'hFF;
            15'd20806: data <= 8'hFF;
            15'd20807: data <= 8'hFF;
            15'd20808: data <= 8'hFF;
            15'd20809: data <= 8'hFF;
            15'd20810: data <= 8'hFF;
            15'd20811: data <= 8'hFF;
            15'd20812: data <= 8'hFF;
            15'd20813: data <= 8'hFF;
            15'd20814: data <= 8'h80;
            15'd20815: data <= 8'h00;
            15'd20816: data <= 8'h00;
            15'd20817: data <= 8'h00;
            15'd20818: data <= 8'h00;
            15'd20819: data <= 8'h00;
            15'd20820: data <= 8'h00;
            15'd20821: data <= 8'h00;
            15'd20822: data <= 8'h00;
            15'd20823: data <= 8'h00;
            15'd20824: data <= 8'h00;
            15'd20825: data <= 8'h03;
            15'd20826: data <= 8'hFF;
            15'd20827: data <= 8'hFF;
            15'd20828: data <= 8'hFF;
            15'd20829: data <= 8'hFF;
            15'd20830: data <= 8'hFF;
            15'd20831: data <= 8'hFF;
            15'd20832: data <= 8'hFF;
            15'd20833: data <= 8'hFF;
            15'd20834: data <= 8'hFF;
            15'd20835: data <= 8'hFF;
            15'd20836: data <= 8'hFF;
            15'd20837: data <= 8'hFF;
            15'd20838: data <= 8'hFF;
            15'd20839: data <= 8'hFF;
            15'd20840: data <= 8'hFF;
            15'd20841: data <= 8'hFF;
            15'd20842: data <= 8'hFF;
            15'd20843: data <= 8'hFF;
            15'd20844: data <= 8'h80;
            15'd20845: data <= 8'h00;
            15'd20846: data <= 8'h00;
            15'd20847: data <= 8'h00;
            15'd20848: data <= 8'h00;
            15'd20849: data <= 8'h00;
            15'd20850: data <= 8'h00;
            15'd20851: data <= 8'h00;
            15'd20852: data <= 8'h00;
            15'd20853: data <= 8'h00;
            15'd20854: data <= 8'h00;
            15'd20855: data <= 8'h03;
            15'd20856: data <= 8'hFF;
            15'd20857: data <= 8'hFF;
            15'd20858: data <= 8'hFF;
            15'd20859: data <= 8'hFF;
            15'd20860: data <= 8'hFF;
            15'd20861: data <= 8'hFF;
            15'd20862: data <= 8'hFF;
            15'd20863: data <= 8'hFF;
            15'd20864: data <= 8'hFF;
            15'd20865: data <= 8'hFF;
            15'd20866: data <= 8'hFF;
            15'd20867: data <= 8'hFF;
            15'd20868: data <= 8'h8F;
            15'd20869: data <= 8'hFF;
            15'd20870: data <= 8'hFF;
            15'd20871: data <= 8'hFF;
            15'd20872: data <= 8'hFF;
            15'd20873: data <= 8'hFF;
            15'd20874: data <= 8'h80;
            15'd20875: data <= 8'h00;
            15'd20876: data <= 8'h00;
            15'd20877: data <= 8'h00;
            15'd20878: data <= 8'h00;
            15'd20879: data <= 8'h00;
            15'd20880: data <= 8'h00;
            15'd20881: data <= 8'h00;
            15'd20882: data <= 8'h00;
            15'd20883: data <= 8'h00;
            15'd20884: data <= 8'h00;
            15'd20885: data <= 8'h03;
            15'd20886: data <= 8'hFF;
            15'd20887: data <= 8'hFF;
            15'd20888: data <= 8'hFF;
            15'd20889: data <= 8'hFF;
            15'd20890: data <= 8'hFB;
            15'd20891: data <= 8'hFF;
            15'd20892: data <= 8'hFF;
            15'd20893: data <= 8'hFF;
            15'd20894: data <= 8'hFE;
            15'd20895: data <= 8'hFF;
            15'd20896: data <= 8'hFF;
            15'd20897: data <= 8'hF8;
            15'd20898: data <= 8'h07;
            15'd20899: data <= 8'hFF;
            15'd20900: data <= 8'hFF;
            15'd20901: data <= 8'hFF;
            15'd20902: data <= 8'hFF;
            15'd20903: data <= 8'hFF;
            15'd20904: data <= 8'h80;
            15'd20905: data <= 8'h00;
            15'd20906: data <= 8'h00;
            15'd20907: data <= 8'h00;
            15'd20908: data <= 8'h00;
            15'd20909: data <= 8'h00;
            15'd20910: data <= 8'h00;
            15'd20911: data <= 8'h00;
            15'd20912: data <= 8'h00;
            15'd20913: data <= 8'h00;
            15'd20914: data <= 8'h00;
            15'd20915: data <= 8'h03;
            15'd20916: data <= 8'hFF;
            15'd20917: data <= 8'hE0;
            15'd20918: data <= 8'h00;
            15'd20919: data <= 8'h3C;
            15'd20920: data <= 8'h0B;
            15'd20921: data <= 8'h7F;
            15'd20922: data <= 8'hFF;
            15'd20923: data <= 8'hFF;
            15'd20924: data <= 8'hFC;
            15'd20925: data <= 8'h7F;
            15'd20926: data <= 8'hFF;
            15'd20927: data <= 8'hC3;
            15'd20928: data <= 8'hF1;
            15'd20929: data <= 8'hFF;
            15'd20930: data <= 8'hFF;
            15'd20931: data <= 8'hE0;
            15'd20932: data <= 8'h1F;
            15'd20933: data <= 8'hFF;
            15'd20934: data <= 8'h80;
            15'd20935: data <= 8'h00;
            15'd20936: data <= 8'h00;
            15'd20937: data <= 8'h00;
            15'd20938: data <= 8'h00;
            15'd20939: data <= 8'h00;
            15'd20940: data <= 8'h00;
            15'd20941: data <= 8'h00;
            15'd20942: data <= 8'h00;
            15'd20943: data <= 8'h00;
            15'd20944: data <= 8'h00;
            15'd20945: data <= 8'h03;
            15'd20946: data <= 8'hFF;
            15'd20947: data <= 8'hFF;
            15'd20948: data <= 8'h77;
            15'd20949: data <= 8'hF0;
            15'd20950: data <= 8'h7B;
            15'd20951: data <= 8'h1F;
            15'd20952: data <= 8'hFF;
            15'd20953: data <= 8'hFE;
            15'd20954: data <= 8'h00;
            15'd20955: data <= 8'h00;
            15'd20956: data <= 8'hFF;
            15'd20957: data <= 8'h9F;
            15'd20958: data <= 8'hFC;
            15'd20959: data <= 8'h3F;
            15'd20960: data <= 8'hF8;
            15'd20961: data <= 8'h7F;
            15'd20962: data <= 8'h9F;
            15'd20963: data <= 8'hFF;
            15'd20964: data <= 8'h80;
            15'd20965: data <= 8'h00;
            15'd20966: data <= 8'h00;
            15'd20967: data <= 8'h00;
            15'd20968: data <= 8'h00;
            15'd20969: data <= 8'h00;
            15'd20970: data <= 8'h00;
            15'd20971: data <= 8'h00;
            15'd20972: data <= 8'h00;
            15'd20973: data <= 8'h00;
            15'd20974: data <= 8'h00;
            15'd20975: data <= 8'h03;
            15'd20976: data <= 8'hFF;
            15'd20977: data <= 8'hFF;
            15'd20978: data <= 8'h77;
            15'd20979: data <= 8'hFE;
            15'd20980: data <= 8'h7B;
            15'd20981: data <= 8'hDF;
            15'd20982: data <= 8'hFF;
            15'd20983: data <= 8'hFF;
            15'd20984: data <= 8'hFE;
            15'd20985: data <= 8'hFF;
            15'd20986: data <= 8'hFF;
            15'd20987: data <= 8'h3F;
            15'd20988: data <= 8'hFF;
            15'd20989: data <= 8'h9F;
            15'd20990: data <= 8'hFB;
            15'd20991: data <= 8'h37;
            15'd20992: data <= 8'h9F;
            15'd20993: data <= 8'hFF;
            15'd20994: data <= 8'h80;
            15'd20995: data <= 8'h00;
            15'd20996: data <= 8'h00;
            15'd20997: data <= 8'h00;
            15'd20998: data <= 8'h00;
            15'd20999: data <= 8'h00;
            15'd21000: data <= 8'h00;
            15'd21001: data <= 8'h00;
            15'd21002: data <= 8'h00;
            15'd21003: data <= 8'h00;
            15'd21004: data <= 8'h00;
            15'd21005: data <= 8'h03;
            15'd21006: data <= 8'hFF;
            15'd21007: data <= 8'hF0;
            15'd21008: data <= 8'h00;
            15'd21009: data <= 8'h3E;
            15'd21010: data <= 8'h7B;
            15'd21011: data <= 8'hFF;
            15'd21012: data <= 8'hFF;
            15'd21013: data <= 8'hFF;
            15'd21014: data <= 8'hC0;
            15'd21015: data <= 8'h0F;
            15'd21016: data <= 8'hFE;
            15'd21017: data <= 8'h7F;
            15'd21018: data <= 8'hFF;
            15'd21019: data <= 8'h9F;
            15'd21020: data <= 8'hFB;
            15'd21021: data <= 8'h37;
            15'd21022: data <= 8'h9F;
            15'd21023: data <= 8'hFF;
            15'd21024: data <= 8'h80;
            15'd21025: data <= 8'h00;
            15'd21026: data <= 8'h00;
            15'd21027: data <= 8'h00;
            15'd21028: data <= 8'h00;
            15'd21029: data <= 8'h00;
            15'd21030: data <= 8'h00;
            15'd21031: data <= 8'h00;
            15'd21032: data <= 8'h00;
            15'd21033: data <= 8'h00;
            15'd21034: data <= 8'h00;
            15'd21035: data <= 8'h03;
            15'd21036: data <= 8'hFF;
            15'd21037: data <= 8'hE7;
            15'd21038: data <= 8'h77;
            15'd21039: data <= 8'h30;
            15'd21040: data <= 8'h00;
            15'd21041: data <= 8'h0F;
            15'd21042: data <= 8'hFF;
            15'd21043: data <= 8'hFF;
            15'd21044: data <= 8'h80;
            15'd21045: data <= 8'h03;
            15'd21046: data <= 8'hFE;
            15'd21047: data <= 8'hEF;
            15'd21048: data <= 8'hFF;
            15'd21049: data <= 8'hDF;
            15'd21050: data <= 8'hFB;
            15'd21051: data <= 8'h27;
            15'd21052: data <= 8'h9F;
            15'd21053: data <= 8'hFF;
            15'd21054: data <= 8'h80;
            15'd21055: data <= 8'h00;
            15'd21056: data <= 8'h00;
            15'd21057: data <= 8'h00;
            15'd21058: data <= 8'h00;
            15'd21059: data <= 8'h00;
            15'd21060: data <= 8'h00;
            15'd21061: data <= 8'h00;
            15'd21062: data <= 8'h00;
            15'd21063: data <= 8'h00;
            15'd21064: data <= 8'h00;
            15'd21065: data <= 8'h03;
            15'd21066: data <= 8'hFF;
            15'd21067: data <= 8'hE7;
            15'd21068: data <= 8'h77;
            15'd21069: data <= 8'h30;
            15'd21070: data <= 8'h00;
            15'd21071: data <= 8'h07;
            15'd21072: data <= 8'hFF;
            15'd21073: data <= 8'hFF;
            15'd21074: data <= 8'h9F;
            15'd21075: data <= 8'hF3;
            15'd21076: data <= 8'hFE;
            15'd21077: data <= 8'hFF;
            15'd21078: data <= 8'hFF;
            15'd21079: data <= 8'hCF;
            15'd21080: data <= 8'hFB;
            15'd21081: data <= 8'h27;
            15'd21082: data <= 8'hBF;
            15'd21083: data <= 8'hFF;
            15'd21084: data <= 8'h80;
            15'd21085: data <= 8'h00;
            15'd21086: data <= 8'h00;
            15'd21087: data <= 8'h00;
            15'd21088: data <= 8'h00;
            15'd21089: data <= 8'h00;
            15'd21090: data <= 8'h00;
            15'd21091: data <= 8'h00;
            15'd21092: data <= 8'h00;
            15'd21093: data <= 8'h00;
            15'd21094: data <= 8'h00;
            15'd21095: data <= 8'h03;
            15'd21096: data <= 8'hFF;
            15'd21097: data <= 8'hE0;
            15'd21098: data <= 8'h00;
            15'd21099: data <= 8'h3E;
            15'd21100: data <= 8'h79;
            15'd21101: data <= 8'hFC;
            15'd21102: data <= 8'h00;
            15'd21103: data <= 8'h03;
            15'd21104: data <= 8'h80;
            15'd21105: data <= 8'h03;
            15'd21106: data <= 8'hFE;
            15'd21107: data <= 8'hFF;
            15'd21108: data <= 8'hFF;
            15'd21109: data <= 8'hE7;
            15'd21110: data <= 8'hFB;
            15'd21111: data <= 8'h27;
            15'd21112: data <= 8'hBF;
            15'd21113: data <= 8'hFF;
            15'd21114: data <= 8'h80;
            15'd21115: data <= 8'h00;
            15'd21116: data <= 8'h00;
            15'd21117: data <= 8'h00;
            15'd21118: data <= 8'h00;
            15'd21119: data <= 8'h00;
            15'd21120: data <= 8'h00;
            15'd21121: data <= 8'h00;
            15'd21122: data <= 8'h00;
            15'd21123: data <= 8'h00;
            15'd21124: data <= 8'h00;
            15'd21125: data <= 8'h03;
            15'd21126: data <= 8'hFF;
            15'd21127: data <= 8'hF7;
            15'd21128: data <= 8'h7F;
            15'd21129: data <= 8'h3E;
            15'd21130: data <= 8'h79;
            15'd21131: data <= 8'hC8;
            15'd21132: data <= 8'h00;
            15'd21133: data <= 8'h03;
            15'd21134: data <= 8'h9F;
            15'd21135: data <= 8'hF3;
            15'd21136: data <= 8'hFE;
            15'd21137: data <= 8'hE3;
            15'd21138: data <= 8'hFF;
            15'd21139: data <= 8'hF7;
            15'd21140: data <= 8'hFB;
            15'd21141: data <= 8'h20;
            15'd21142: data <= 8'h0F;
            15'd21143: data <= 8'hFF;
            15'd21144: data <= 8'h80;
            15'd21145: data <= 8'h00;
            15'd21146: data <= 8'h00;
            15'd21147: data <= 8'h00;
            15'd21148: data <= 8'h00;
            15'd21149: data <= 8'h00;
            15'd21150: data <= 8'h00;
            15'd21151: data <= 8'h00;
            15'd21152: data <= 8'h00;
            15'd21153: data <= 8'h00;
            15'd21154: data <= 8'h00;
            15'd21155: data <= 8'h03;
            15'd21156: data <= 8'hFF;
            15'd21157: data <= 8'hFF;
            15'd21158: data <= 8'h7F;
            15'd21159: data <= 8'hFE;
            15'd21160: data <= 8'h0D;
            15'd21161: data <= 8'h9F;
            15'd21162: data <= 8'hFF;
            15'd21163: data <= 8'hFF;
            15'd21164: data <= 8'h9F;
            15'd21165: data <= 8'hF3;
            15'd21166: data <= 8'hFE;
            15'd21167: data <= 8'h05;
            15'd21168: data <= 8'hFF;
            15'd21169: data <= 8'hF3;
            15'd21170: data <= 8'hFB;
            15'd21171: data <= 8'h3F;
            15'd21172: data <= 8'hEF;
            15'd21173: data <= 8'hFF;
            15'd21174: data <= 8'h80;
            15'd21175: data <= 8'h00;
            15'd21176: data <= 8'h00;
            15'd21177: data <= 8'h00;
            15'd21178: data <= 8'h00;
            15'd21179: data <= 8'h00;
            15'd21180: data <= 8'h00;
            15'd21181: data <= 8'h00;
            15'd21182: data <= 8'h00;
            15'd21183: data <= 8'h00;
            15'd21184: data <= 8'h00;
            15'd21185: data <= 8'h03;
            15'd21186: data <= 8'hFF;
            15'd21187: data <= 8'hC0;
            15'd21188: data <= 8'h00;
            15'd21189: data <= 8'h10;
            15'd21190: data <= 8'h1D;
            15'd21191: data <= 8'h3F;
            15'd21192: data <= 8'hFF;
            15'd21193: data <= 8'hFF;
            15'd21194: data <= 8'h80;
            15'd21195: data <= 8'h03;
            15'd21196: data <= 8'hFF;
            15'd21197: data <= 8'h01;
            15'd21198: data <= 8'hFF;
            15'd21199: data <= 8'hFB;
            15'd21200: data <= 8'hFB;
            15'd21201: data <= 8'h3F;
            15'd21202: data <= 8'hEF;
            15'd21203: data <= 8'hFF;
            15'd21204: data <= 8'h80;
            15'd21205: data <= 8'h00;
            15'd21206: data <= 8'h00;
            15'd21207: data <= 8'h00;
            15'd21208: data <= 8'h00;
            15'd21209: data <= 8'h00;
            15'd21210: data <= 8'h00;
            15'd21211: data <= 8'h00;
            15'd21212: data <= 8'h00;
            15'd21213: data <= 8'h00;
            15'd21214: data <= 8'h00;
            15'd21215: data <= 8'h03;
            15'd21216: data <= 8'hFF;
            15'd21217: data <= 8'hFC;
            15'd21218: data <= 8'hF9;
            15'd21219: data <= 8'hF2;
            15'd21220: data <= 8'h7C;
            15'd21221: data <= 8'h7F;
            15'd21222: data <= 8'hFF;
            15'd21223: data <= 8'hFF;
            15'd21224: data <= 8'h9F;
            15'd21225: data <= 8'hF3;
            15'd21226: data <= 8'hFF;
            15'd21227: data <= 8'h9F;
            15'd21228: data <= 8'hFF;
            15'd21229: data <= 8'hFB;
            15'd21230: data <= 8'hFB;
            15'd21231: data <= 8'h3F;
            15'd21232: data <= 8'hEF;
            15'd21233: data <= 8'hFF;
            15'd21234: data <= 8'h80;
            15'd21235: data <= 8'h00;
            15'd21236: data <= 8'h00;
            15'd21237: data <= 8'h00;
            15'd21238: data <= 8'h00;
            15'd21239: data <= 8'h00;
            15'd21240: data <= 8'h00;
            15'd21241: data <= 8'h00;
            15'd21242: data <= 8'h00;
            15'd21243: data <= 8'h00;
            15'd21244: data <= 8'h00;
            15'd21245: data <= 8'h03;
            15'd21246: data <= 8'hFF;
            15'd21247: data <= 8'hFD;
            15'd21248: data <= 8'hFB;
            15'd21249: data <= 8'hFE;
            15'd21250: data <= 8'h7C;
            15'd21251: data <= 8'hFF;
            15'd21252: data <= 8'hFF;
            15'd21253: data <= 8'hFF;
            15'd21254: data <= 8'h80;
            15'd21255: data <= 8'h03;
            15'd21256: data <= 8'hFF;
            15'd21257: data <= 8'hAD;
            15'd21258: data <= 8'hFF;
            15'd21259: data <= 8'hF9;
            15'd21260: data <= 8'hF8;
            15'd21261: data <= 8'h00;
            15'd21262: data <= 8'h2F;
            15'd21263: data <= 8'hFF;
            15'd21264: data <= 8'h80;
            15'd21265: data <= 8'h00;
            15'd21266: data <= 8'h00;
            15'd21267: data <= 8'h00;
            15'd21268: data <= 8'h00;
            15'd21269: data <= 8'h00;
            15'd21270: data <= 8'h00;
            15'd21271: data <= 8'h00;
            15'd21272: data <= 8'h00;
            15'd21273: data <= 8'h00;
            15'd21274: data <= 8'h00;
            15'd21275: data <= 8'h03;
            15'd21276: data <= 8'hFF;
            15'd21277: data <= 8'hFC;
            15'd21278: data <= 8'h27;
            15'd21279: data <= 8'hFE;
            15'd21280: data <= 8'h70;
            15'd21281: data <= 8'hE7;
            15'd21282: data <= 8'hFF;
            15'd21283: data <= 8'hFF;
            15'd21284: data <= 8'h80;
            15'd21285: data <= 8'h03;
            15'd21286: data <= 8'hFF;
            15'd21287: data <= 8'hAE;
            15'd21288: data <= 8'h67;
            15'd21289: data <= 8'hFD;
            15'd21290: data <= 8'hFB;
            15'd21291: data <= 8'h3F;
            15'd21292: data <= 8'hEF;
            15'd21293: data <= 8'hFF;
            15'd21294: data <= 8'h80;
            15'd21295: data <= 8'h00;
            15'd21296: data <= 8'h00;
            15'd21297: data <= 8'h00;
            15'd21298: data <= 8'h00;
            15'd21299: data <= 8'h00;
            15'd21300: data <= 8'h00;
            15'd21301: data <= 8'h00;
            15'd21302: data <= 8'h00;
            15'd21303: data <= 8'h00;
            15'd21304: data <= 8'h00;
            15'd21305: data <= 8'h03;
            15'd21306: data <= 8'hFF;
            15'd21307: data <= 8'hFF;
            15'd21308: data <= 8'h87;
            15'd21309: data <= 8'hFE;
            15'd21310: data <= 8'h66;
            15'd21311: data <= 8'h6F;
            15'd21312: data <= 8'hFF;
            15'd21313: data <= 8'hFF;
            15'd21314: data <= 8'h9F;
            15'd21315: data <= 8'hF3;
            15'd21316: data <= 8'hFF;
            15'd21317: data <= 8'hB7;
            15'd21318: data <= 8'h8F;
            15'd21319: data <= 8'hFC;
            15'd21320: data <= 8'hFF;
            15'd21321: data <= 8'hFF;
            15'd21322: data <= 8'hEF;
            15'd21323: data <= 8'hFF;
            15'd21324: data <= 8'h80;
            15'd21325: data <= 8'h00;
            15'd21326: data <= 8'h00;
            15'd21327: data <= 8'h00;
            15'd21328: data <= 8'h00;
            15'd21329: data <= 8'h00;
            15'd21330: data <= 8'h00;
            15'd21331: data <= 8'h00;
            15'd21332: data <= 8'h00;
            15'd21333: data <= 8'h00;
            15'd21334: data <= 8'h00;
            15'd21335: data <= 8'h03;
            15'd21336: data <= 8'hFF;
            15'd21337: data <= 8'hFC;
            15'd21338: data <= 8'h30;
            15'd21339: data <= 8'h7E;
            15'd21340: data <= 8'h4F;
            15'd21341: data <= 8'h2F;
            15'd21342: data <= 8'hFF;
            15'd21343: data <= 8'hFE;
            15'd21344: data <= 8'h00;
            15'd21345: data <= 8'h00;
            15'd21346: data <= 8'hFF;
            15'd21347: data <= 8'hF7;
            15'd21348: data <= 8'hFF;
            15'd21349: data <= 8'hFC;
            15'd21350: data <= 8'hFF;
            15'd21351: data <= 8'hFC;
            15'd21352: data <= 8'h0F;
            15'd21353: data <= 8'hFF;
            15'd21354: data <= 8'h80;
            15'd21355: data <= 8'h00;
            15'd21356: data <= 8'h00;
            15'd21357: data <= 8'h00;
            15'd21358: data <= 8'h00;
            15'd21359: data <= 8'h00;
            15'd21360: data <= 8'h00;
            15'd21361: data <= 8'h00;
            15'd21362: data <= 8'h00;
            15'd21363: data <= 8'h00;
            15'd21364: data <= 8'h00;
            15'd21365: data <= 8'h03;
            15'd21366: data <= 8'hFF;
            15'd21367: data <= 8'hE1;
            15'd21368: data <= 8'hFE;
            15'd21369: data <= 8'h38;
            15'd21370: data <= 8'hFF;
            15'd21371: data <= 8'h8F;
            15'd21372: data <= 8'hFF;
            15'd21373: data <= 8'hFE;
            15'd21374: data <= 8'h00;
            15'd21375: data <= 8'h00;
            15'd21376: data <= 8'hFF;
            15'd21377: data <= 8'hFB;
            15'd21378: data <= 8'hFF;
            15'd21379: data <= 8'hFE;
            15'd21380: data <= 8'hFF;
            15'd21381: data <= 8'hFC;
            15'd21382: data <= 8'h1F;
            15'd21383: data <= 8'hFF;
            15'd21384: data <= 8'h80;
            15'd21385: data <= 8'h00;
            15'd21386: data <= 8'h00;
            15'd21387: data <= 8'h00;
            15'd21388: data <= 8'h00;
            15'd21389: data <= 8'h00;
            15'd21390: data <= 8'h00;
            15'd21391: data <= 8'h00;
            15'd21392: data <= 8'h00;
            15'd21393: data <= 8'h00;
            15'd21394: data <= 8'h00;
            15'd21395: data <= 8'h03;
            15'd21396: data <= 8'hFF;
            15'd21397: data <= 8'hFF;
            15'd21398: data <= 8'hFF;
            15'd21399: data <= 8'hFF;
            15'd21400: data <= 8'hFF;
            15'd21401: data <= 8'hFF;
            15'd21402: data <= 8'hFF;
            15'd21403: data <= 8'hFF;
            15'd21404: data <= 8'hFF;
            15'd21405: data <= 8'hFF;
            15'd21406: data <= 8'hFF;
            15'd21407: data <= 8'hBD;
            15'd21408: data <= 8'hFF;
            15'd21409: data <= 8'hFE;
            15'd21410: data <= 8'hFF;
            15'd21411: data <= 8'hFF;
            15'd21412: data <= 8'hFF;
            15'd21413: data <= 8'hFF;
            15'd21414: data <= 8'h80;
            15'd21415: data <= 8'h00;
            15'd21416: data <= 8'h00;
            15'd21417: data <= 8'h00;
            15'd21418: data <= 8'h00;
            15'd21419: data <= 8'h00;
            15'd21420: data <= 8'h00;
            15'd21421: data <= 8'h00;
            15'd21422: data <= 8'h00;
            15'd21423: data <= 8'h00;
            15'd21424: data <= 8'h00;
            15'd21425: data <= 8'h03;
            15'd21426: data <= 8'hFF;
            15'd21427: data <= 8'hFF;
            15'd21428: data <= 8'hFF;
            15'd21429: data <= 8'hFF;
            15'd21430: data <= 8'hFF;
            15'd21431: data <= 8'hFF;
            15'd21432: data <= 8'hFF;
            15'd21433: data <= 8'hFF;
            15'd21434: data <= 8'hFF;
            15'd21435: data <= 8'hFF;
            15'd21436: data <= 8'hFF;
            15'd21437: data <= 8'hBE;
            15'd21438: data <= 8'h7F;
            15'd21439: data <= 8'hFE;
            15'd21440: data <= 8'h7F;
            15'd21441: data <= 8'hFF;
            15'd21442: data <= 8'hFF;
            15'd21443: data <= 8'hFF;
            15'd21444: data <= 8'h80;
            15'd21445: data <= 8'h00;
            15'd21446: data <= 8'h00;
            15'd21447: data <= 8'h00;
            15'd21448: data <= 8'h00;
            15'd21449: data <= 8'h00;
            15'd21450: data <= 8'h00;
            15'd21451: data <= 8'h00;
            15'd21452: data <= 8'h00;
            15'd21453: data <= 8'h00;
            15'd21454: data <= 8'h00;
            15'd21455: data <= 8'h03;
            15'd21456: data <= 8'hFF;
            15'd21457: data <= 8'hFF;
            15'd21458: data <= 8'hFF;
            15'd21459: data <= 8'hFF;
            15'd21460: data <= 8'hFF;
            15'd21461: data <= 8'hFF;
            15'd21462: data <= 8'hFF;
            15'd21463: data <= 8'hFF;
            15'd21464: data <= 8'hFF;
            15'd21465: data <= 8'hFF;
            15'd21466: data <= 8'hFF;
            15'd21467: data <= 8'hBF;
            15'd21468: data <= 8'h03;
            15'd21469: data <= 8'hFE;
            15'd21470: data <= 8'h7F;
            15'd21471: data <= 8'hFF;
            15'd21472: data <= 8'hFF;
            15'd21473: data <= 8'hFF;
            15'd21474: data <= 8'h80;
            15'd21475: data <= 8'h00;
            15'd21476: data <= 8'h00;
            15'd21477: data <= 8'h00;
            15'd21478: data <= 8'h00;
            15'd21479: data <= 8'h00;
            15'd21480: data <= 8'h00;
            15'd21481: data <= 8'h00;
            15'd21482: data <= 8'h00;
            15'd21483: data <= 8'h00;
            15'd21484: data <= 8'h00;
            15'd21485: data <= 8'h03;
            15'd21486: data <= 8'hFF;
            15'd21487: data <= 8'hFF;
            15'd21488: data <= 8'hFF;
            15'd21489: data <= 8'hFF;
            15'd21490: data <= 8'hFF;
            15'd21491: data <= 8'hFF;
            15'd21492: data <= 8'hFF;
            15'd21493: data <= 8'hFF;
            15'd21494: data <= 8'hFF;
            15'd21495: data <= 8'hFF;
            15'd21496: data <= 8'hFF;
            15'd21497: data <= 8'hBF;
            15'd21498: data <= 8'hFF;
            15'd21499: data <= 8'hFF;
            15'd21500: data <= 8'h7F;
            15'd21501: data <= 8'hFF;
            15'd21502: data <= 8'hFF;
            15'd21503: data <= 8'hFF;
            15'd21504: data <= 8'h80;
            15'd21505: data <= 8'h00;
            15'd21506: data <= 8'h00;
            15'd21507: data <= 8'h00;
            15'd21508: data <= 8'h00;
            15'd21509: data <= 8'h00;
            15'd21510: data <= 8'h00;
            15'd21511: data <= 8'h00;
            15'd21512: data <= 8'h00;
            15'd21513: data <= 8'h00;
            15'd21514: data <= 8'h00;
            15'd21515: data <= 8'h03;
            15'd21516: data <= 8'hFF;
            15'd21517: data <= 8'hFF;
            15'd21518: data <= 8'hFF;
            15'd21519: data <= 8'hFF;
            15'd21520: data <= 8'hFF;
            15'd21521: data <= 8'hFF;
            15'd21522: data <= 8'hFF;
            15'd21523: data <= 8'hFF;
            15'd21524: data <= 8'hFF;
            15'd21525: data <= 8'hFF;
            15'd21526: data <= 8'hFF;
            15'd21527: data <= 8'hBF;
            15'd21528: data <= 8'hFF;
            15'd21529: data <= 8'hFF;
            15'd21530: data <= 8'h7F;
            15'd21531: data <= 8'hFF;
            15'd21532: data <= 8'hFF;
            15'd21533: data <= 8'hFF;
            15'd21534: data <= 8'h80;
            15'd21535: data <= 8'h00;
            15'd21536: data <= 8'h00;
            15'd21537: data <= 8'h00;
            15'd21538: data <= 8'h00;
            15'd21539: data <= 8'h00;
            15'd21540: data <= 8'h00;
            15'd21541: data <= 8'h00;
            15'd21542: data <= 8'h00;
            15'd21543: data <= 8'h00;
            15'd21544: data <= 8'h00;
            15'd21545: data <= 8'h03;
            15'd21546: data <= 8'hFF;
            15'd21547: data <= 8'hFF;
            15'd21548: data <= 8'hFF;
            15'd21549: data <= 8'hFF;
            15'd21550: data <= 8'hFF;
            15'd21551: data <= 8'hFF;
            15'd21552: data <= 8'hFF;
            15'd21553: data <= 8'hFF;
            15'd21554: data <= 8'hFF;
            15'd21555: data <= 8'hFF;
            15'd21556: data <= 8'hFF;
            15'd21557: data <= 8'hBF;
            15'd21558: data <= 8'hFF;
            15'd21559: data <= 8'hFF;
            15'd21560: data <= 8'hFF;
            15'd21561: data <= 8'hFF;
            15'd21562: data <= 8'hFF;
            15'd21563: data <= 8'hFF;
            15'd21564: data <= 8'h80;
            15'd21565: data <= 8'h00;
            15'd21566: data <= 8'h00;
            15'd21567: data <= 8'h00;
            15'd21568: data <= 8'h00;
            15'd21569: data <= 8'h00;
            15'd21570: data <= 8'h00;
            15'd21571: data <= 8'h00;
            15'd21572: data <= 8'h00;
            15'd21573: data <= 8'h00;
            15'd21574: data <= 8'h00;
            15'd21575: data <= 8'h03;
            15'd21576: data <= 8'hFF;
            15'd21577: data <= 8'hFF;
            15'd21578: data <= 8'hFF;
            15'd21579: data <= 8'hFF;
            15'd21580: data <= 8'hFF;
            15'd21581: data <= 8'hFF;
            15'd21582: data <= 8'hFF;
            15'd21583: data <= 8'hFF;
            15'd21584: data <= 8'hFF;
            15'd21585: data <= 8'hFF;
            15'd21586: data <= 8'hFF;
            15'd21587: data <= 8'hFF;
            15'd21588: data <= 8'hFF;
            15'd21589: data <= 8'hFF;
            15'd21590: data <= 8'hFF;
            15'd21591: data <= 8'hFF;
            15'd21592: data <= 8'hFF;
            15'd21593: data <= 8'hFF;
            15'd21594: data <= 8'h80;
            15'd21595: data <= 8'h00;
            15'd21596: data <= 8'h00;
            15'd21597: data <= 8'h00;
            15'd21598: data <= 8'h00;
            15'd21599: data <= 8'h00;
            default: data <= 8'h00;
        endcase
    end

endmodule
