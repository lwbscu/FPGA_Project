// tone.v - 音调转换模块
// 将按键信息转换为对应的PWM周期值
// 系统时钟12MHz，根据音调频率计算周期值

module tone(
    input   [15:0]  key_in,     // 按键输入（one-hot编码）
    output reg [15:0] cycle     // PWM周期输出
);

// 组合逻辑：根据按键输入选择对应的周期值
// 周期值 = 12MHz / 音调频率
always @(key_in) begin
    case(key_in)
        16'h0001: cycle = 16'd45872;    // K1  - 低音1 (261.6Hz)
        16'h0002: cycle = 16'd40858;    // K2  - 低音2 (293.7Hz)
        16'h0004: cycle = 16'd36408;    // K3  - 低音3 (329.6Hz)
        16'h0008: cycle = 16'd34364;    // K4  - 低音4 (349.2Hz)
        16'h0010: cycle = 16'd30612;    // K5  - 低音5 (392Hz)
        16'h0020: cycle = 16'd27273;    // K6  - 低音6 (440Hz)
        16'h0040: cycle = 16'd24296;    // K7  - 低音7 (493.9Hz)
        16'h0080: cycle = 16'd22931;    // K8  - 中音1 (523.3Hz)
        16'h0100: cycle = 16'd20432;    // K9  - 中音2 (587.3Hz)
        16'h0200: cycle = 16'd18201;    // K10 - 中音3 (659.3Hz)
        16'h0400: cycle = 16'd17180;    // K11 - 中音4 (698.5Hz)
        16'h0800: cycle = 16'd15306;    // K12 - 中音5 (784Hz)
        16'h1000: cycle = 16'd13636;    // K13 - 中音6 (880Hz)
        16'h2000: cycle = 16'd12148;    // K14 - 中音7 (987.8Hz)
        16'h4000: cycle = 16'd11478;    // K15 - 高音1 (1045.5Hz)
        16'h8000: cycle = 16'd10215;    // K16 - 高音2 (1174.7Hz)
        default:  cycle = 16'd0;         // 无按键按下，输出0（静音）
    endcase
end

endmodule