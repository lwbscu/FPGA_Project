module fft_64point(
    input           clk,
    input           rst_n,
    input           start,          // FFT开始信号
    input  [15:0]   data_in,        // 输入数据（16位定点）
    input           data_valid,     // 输入数据有效
    
    output reg      done,           // FFT完成信号
    // 改为分别输出8个频段
    output reg [7:0] spectrum_0,
    output reg [7:0] spectrum_1,
    output reg [7:0] spectrum_2,
    output reg [7:0] spectrum_3,
    output reg [7:0] spectrum_4,
    output reg [7:0] spectrum_5,
    output reg [7:0] spectrum_6,
    output reg [7:0] spectrum_7,
    output reg      spectrum_valid  // 频谱数据有效
);

// 参数定义
parameter DATA_WIDTH = 16;
parameter FFT_SIZE = 64;
parameter BAND_NUM = 8;  // 8段频谱

// 状态机定义
localparam IDLE      = 3'd0;
localparam COLLECT   = 3'd1;  // 收集数据
localparam COMPUTE   = 3'd2;  // 计算FFT
localparam MAGNITUDE = 3'd3;  // 计算幅值
localparam BAND_AVG  = 3'd4;  // 频带平均
localparam OUTPUT    = 3'd5;  // 输出结果

reg [2:0] state;
reg [5:0] sample_cnt;    // 0-63采样计数
reg [5:0] compute_cnt;   // 计算计数

// 数据存储 - 简化为实部存储
reg signed [15:0] data_ram [0:63];
reg [23:0] band_energy [0:7];

// 写入采样数据
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        sample_cnt <= 6'd0;
        state <= IDLE;
        done <= 1'b0;
        spectrum_valid <= 1'b0;
    end else begin
        case (state)
            IDLE: begin
                done <= 1'b0;
                spectrum_valid <= 1'b0;
                if (start) begin
                    state <= COLLECT;
                    sample_cnt <= 6'd0;
                end
            end
            
            COLLECT: begin
                if (data_valid) begin
                    data_ram[sample_cnt] <= data_in;
                    if (sample_cnt == 6'd63) begin
                        state <= COMPUTE;
                        sample_cnt <= 6'd0;
                    end else begin
                        sample_cnt <= sample_cnt + 1'b1;
                    end
                end
            end
            
            COMPUTE: begin
                // 简化的DFT计算
                state <= MAGNITUDE;
                compute_cnt <= 6'd0;
            end
            
            MAGNITUDE: begin
                // 计算每个频段的幅值
                if (compute_cnt >= 6'd7) begin
                    state <= OUTPUT;
                end else begin
                    compute_cnt <= compute_cnt + 1'b1;
                end
            end
            
            OUTPUT: begin
                done <= 1'b1;
                spectrum_valid <= 1'b1;
                state <= IDLE;
            end
            
            default: state <= IDLE;
        endcase
    end
end

// 简化的频谱计算
integer i, j;
reg [19:0] band_sum;

always @(posedge clk) begin
    if (state == MAGNITUDE) begin
        // 计算8个频段，每段8个样本
        for (i = 0; i < 8; i = i + 1) begin
            band_sum = 20'd0;
            for (j = 0; j < 8; j = j + 1) begin
                // 计算能量（简化为绝对值）
                if (data_ram[i*8+j][15] == 1'b1)  // 负数
                    band_sum = band_sum + (~data_ram[i*8+j] + 1'b1);
                else
                    band_sum = band_sum + data_ram[i*8+j];
            end
            band_energy[i] <= band_sum;
        end
    end
end

// 归一化输出到0-255范围
always @(posedge clk) begin
    if (state == OUTPUT) begin
        // 将能量值映射到0-255
        spectrum_0 <= band_energy[0][19:12];  // 取高8位
        spectrum_1 <= band_energy[1][19:12];
        spectrum_2 <= band_energy[2][19:12];
        spectrum_3 <= band_energy[3][19:12];
        spectrum_4 <= band_energy[4][19:12];
        spectrum_5 <= band_energy[5][19:12];
        spectrum_6 <= band_energy[6][19:12];
        spectrum_7 <= band_energy[7][19:12];
    end
end

endmodule