// �Զ����ɵ�ROMģ��
// ͼƬ�ߴ�: 320 x 240
// ��ɫ��ʽ: �ڰ�(1λ)
// ���ݴ�С: 9600 �ֽ�
// ���ɹ���: image_processor.py

module image_0_rom (
    input wire clk,
    input wire [13:0] addr,
    output reg [7:0] data
);

    // ROM���ݴ洢 (9600 ����ַ)
    always @(posedge clk) begin
        case (addr)
            14'd0: data <= 8'h00;
            14'd1: data <= 8'h00;
            14'd2: data <= 8'h00;
            14'd3: data <= 8'h00;
            14'd4: data <= 8'h00;
            14'd5: data <= 8'h00;
            14'd6: data <= 8'h0F;
            14'd7: data <= 8'hFF;
            14'd8: data <= 8'hFF;
            14'd9: data <= 8'hFF;
            14'd10: data <= 8'hFF;
            14'd11: data <= 8'hFF;
            14'd12: data <= 8'hFF;
            14'd13: data <= 8'hFF;
            14'd14: data <= 8'hFF;
            14'd15: data <= 8'hFF;
            14'd16: data <= 8'hFF;
            14'd17: data <= 8'hFF;
            14'd18: data <= 8'hFF;
            14'd19: data <= 8'hFF;
            14'd20: data <= 8'hFF;
            14'd21: data <= 8'hFF;
            14'd22: data <= 8'hFF;
            14'd23: data <= 8'hFF;
            14'd24: data <= 8'hFF;
            14'd25: data <= 8'hFF;
            14'd26: data <= 8'hFF;
            14'd27: data <= 8'hFF;
            14'd28: data <= 8'hFF;
            14'd29: data <= 8'hFF;
            14'd30: data <= 8'hFF;
            14'd31: data <= 8'hFF;
            14'd32: data <= 8'hFF;
            14'd33: data <= 8'hF0;
            14'd34: data <= 8'h00;
            14'd35: data <= 8'h00;
            14'd36: data <= 8'h00;
            14'd37: data <= 8'h00;
            14'd38: data <= 8'h00;
            14'd39: data <= 8'h00;
            14'd40: data <= 8'h00;
            14'd41: data <= 8'h00;
            14'd42: data <= 8'h00;
            14'd43: data <= 8'h00;
            14'd44: data <= 8'h00;
            14'd45: data <= 8'h00;
            14'd46: data <= 8'h0F;
            14'd47: data <= 8'hFF;
            14'd48: data <= 8'hFF;
            14'd49: data <= 8'hFF;
            14'd50: data <= 8'hFF;
            14'd51: data <= 8'hFF;
            14'd52: data <= 8'hFF;
            14'd53: data <= 8'hFF;
            14'd54: data <= 8'hFF;
            14'd55: data <= 8'hFF;
            14'd56: data <= 8'hFF;
            14'd57: data <= 8'hFF;
            14'd58: data <= 8'hFF;
            14'd59: data <= 8'hFF;
            14'd60: data <= 8'hFF;
            14'd61: data <= 8'hFF;
            14'd62: data <= 8'hFF;
            14'd63: data <= 8'hFF;
            14'd64: data <= 8'hFF;
            14'd65: data <= 8'hFF;
            14'd66: data <= 8'hFF;
            14'd67: data <= 8'hFF;
            14'd68: data <= 8'hFF;
            14'd69: data <= 8'hFF;
            14'd70: data <= 8'hFF;
            14'd71: data <= 8'hFF;
            14'd72: data <= 8'hFF;
            14'd73: data <= 8'hF0;
            14'd74: data <= 8'h00;
            14'd75: data <= 8'h00;
            14'd76: data <= 8'h00;
            14'd77: data <= 8'h00;
            14'd78: data <= 8'h00;
            14'd79: data <= 8'h00;
            14'd80: data <= 8'h00;
            14'd81: data <= 8'h00;
            14'd82: data <= 8'h00;
            14'd83: data <= 8'h00;
            14'd84: data <= 8'h00;
            14'd85: data <= 8'h00;
            14'd86: data <= 8'h0F;
            14'd87: data <= 8'hFF;
            14'd88: data <= 8'hFF;
            14'd89: data <= 8'hFF;
            14'd90: data <= 8'hFF;
            14'd91: data <= 8'hFF;
            14'd92: data <= 8'hFF;
            14'd93: data <= 8'hFF;
            14'd94: data <= 8'hFF;
            14'd95: data <= 8'hFF;
            14'd96: data <= 8'hFF;
            14'd97: data <= 8'hFF;
            14'd98: data <= 8'hFF;
            14'd99: data <= 8'hFF;
            14'd100: data <= 8'hFF;
            14'd101: data <= 8'hFF;
            14'd102: data <= 8'hFF;
            14'd103: data <= 8'hFF;
            14'd104: data <= 8'hFF;
            14'd105: data <= 8'hFF;
            14'd106: data <= 8'hFF;
            14'd107: data <= 8'hFF;
            14'd108: data <= 8'hFF;
            14'd109: data <= 8'hFF;
            14'd110: data <= 8'hFF;
            14'd111: data <= 8'hFF;
            14'd112: data <= 8'hFF;
            14'd113: data <= 8'hF0;
            14'd114: data <= 8'h00;
            14'd115: data <= 8'h00;
            14'd116: data <= 8'h00;
            14'd117: data <= 8'h00;
            14'd118: data <= 8'h00;
            14'd119: data <= 8'h00;
            14'd120: data <= 8'h00;
            14'd121: data <= 8'h00;
            14'd122: data <= 8'h00;
            14'd123: data <= 8'h00;
            14'd124: data <= 8'h00;
            14'd125: data <= 8'h00;
            14'd126: data <= 8'h0F;
            14'd127: data <= 8'hFF;
            14'd128: data <= 8'hFF;
            14'd129: data <= 8'hFF;
            14'd130: data <= 8'hFF;
            14'd131: data <= 8'hFF;
            14'd132: data <= 8'hFF;
            14'd133: data <= 8'hFF;
            14'd134: data <= 8'hFF;
            14'd135: data <= 8'hFF;
            14'd136: data <= 8'hFF;
            14'd137: data <= 8'hFF;
            14'd138: data <= 8'hFF;
            14'd139: data <= 8'hFF;
            14'd140: data <= 8'hFF;
            14'd141: data <= 8'hFF;
            14'd142: data <= 8'hFF;
            14'd143: data <= 8'hFF;
            14'd144: data <= 8'hFF;
            14'd145: data <= 8'hFF;
            14'd146: data <= 8'hFF;
            14'd147: data <= 8'hFF;
            14'd148: data <= 8'hFF;
            14'd149: data <= 8'hFF;
            14'd150: data <= 8'hFF;
            14'd151: data <= 8'hFF;
            14'd152: data <= 8'hFF;
            14'd153: data <= 8'hF0;
            14'd154: data <= 8'h00;
            14'd155: data <= 8'h00;
            14'd156: data <= 8'h00;
            14'd157: data <= 8'h00;
            14'd158: data <= 8'h00;
            14'd159: data <= 8'h00;
            14'd160: data <= 8'h00;
            14'd161: data <= 8'h00;
            14'd162: data <= 8'h00;
            14'd163: data <= 8'h00;
            14'd164: data <= 8'h00;
            14'd165: data <= 8'h00;
            14'd166: data <= 8'h0F;
            14'd167: data <= 8'hFF;
            14'd168: data <= 8'hFF;
            14'd169: data <= 8'hFF;
            14'd170: data <= 8'hFF;
            14'd171: data <= 8'hFF;
            14'd172: data <= 8'hFF;
            14'd173: data <= 8'hFF;
            14'd174: data <= 8'hFF;
            14'd175: data <= 8'hFF;
            14'd176: data <= 8'hFF;
            14'd177: data <= 8'hFF;
            14'd178: data <= 8'hFF;
            14'd179: data <= 8'hFF;
            14'd180: data <= 8'hFF;
            14'd181: data <= 8'hFF;
            14'd182: data <= 8'hFF;
            14'd183: data <= 8'hFF;
            14'd184: data <= 8'hFF;
            14'd185: data <= 8'hFF;
            14'd186: data <= 8'hFF;
            14'd187: data <= 8'hFF;
            14'd188: data <= 8'hFF;
            14'd189: data <= 8'hFF;
            14'd190: data <= 8'hFF;
            14'd191: data <= 8'hFF;
            14'd192: data <= 8'hFF;
            14'd193: data <= 8'hF0;
            14'd194: data <= 8'h00;
            14'd195: data <= 8'h00;
            14'd196: data <= 8'h00;
            14'd197: data <= 8'h00;
            14'd198: data <= 8'h00;
            14'd199: data <= 8'h00;
            14'd200: data <= 8'h00;
            14'd201: data <= 8'h00;
            14'd202: data <= 8'h00;
            14'd203: data <= 8'h00;
            14'd204: data <= 8'h00;
            14'd205: data <= 8'h00;
            14'd206: data <= 8'h0F;
            14'd207: data <= 8'hFF;
            14'd208: data <= 8'hFF;
            14'd209: data <= 8'hFF;
            14'd210: data <= 8'hFF;
            14'd211: data <= 8'hFF;
            14'd212: data <= 8'hFF;
            14'd213: data <= 8'hFF;
            14'd214: data <= 8'hFF;
            14'd215: data <= 8'hFF;
            14'd216: data <= 8'hFF;
            14'd217: data <= 8'hFF;
            14'd218: data <= 8'hFF;
            14'd219: data <= 8'hFF;
            14'd220: data <= 8'hFF;
            14'd221: data <= 8'hFF;
            14'd222: data <= 8'hFF;
            14'd223: data <= 8'hFF;
            14'd224: data <= 8'hFF;
            14'd225: data <= 8'hFF;
            14'd226: data <= 8'hFF;
            14'd227: data <= 8'hFF;
            14'd228: data <= 8'hFF;
            14'd229: data <= 8'hFF;
            14'd230: data <= 8'hFF;
            14'd231: data <= 8'hFF;
            14'd232: data <= 8'hFF;
            14'd233: data <= 8'hF0;
            14'd234: data <= 8'h00;
            14'd235: data <= 8'h00;
            14'd236: data <= 8'h00;
            14'd237: data <= 8'h00;
            14'd238: data <= 8'h00;
            14'd239: data <= 8'h00;
            14'd240: data <= 8'h00;
            14'd241: data <= 8'h00;
            14'd242: data <= 8'h00;
            14'd243: data <= 8'h00;
            14'd244: data <= 8'h00;
            14'd245: data <= 8'h00;
            14'd246: data <= 8'h0F;
            14'd247: data <= 8'hFF;
            14'd248: data <= 8'hFF;
            14'd249: data <= 8'hFF;
            14'd250: data <= 8'hFF;
            14'd251: data <= 8'hFF;
            14'd252: data <= 8'hFF;
            14'd253: data <= 8'hFF;
            14'd254: data <= 8'hFF;
            14'd255: data <= 8'hFF;
            14'd256: data <= 8'hFF;
            14'd257: data <= 8'hFF;
            14'd258: data <= 8'hFF;
            14'd259: data <= 8'hFF;
            14'd260: data <= 8'hFF;
            14'd261: data <= 8'hFF;
            14'd262: data <= 8'hFF;
            14'd263: data <= 8'hFF;
            14'd264: data <= 8'hFF;
            14'd265: data <= 8'hFF;
            14'd266: data <= 8'hFF;
            14'd267: data <= 8'hFF;
            14'd268: data <= 8'hFF;
            14'd269: data <= 8'hFF;
            14'd270: data <= 8'hFF;
            14'd271: data <= 8'hFF;
            14'd272: data <= 8'hFF;
            14'd273: data <= 8'hF0;
            14'd274: data <= 8'h00;
            14'd275: data <= 8'h00;
            14'd276: data <= 8'h00;
            14'd277: data <= 8'h00;
            14'd278: data <= 8'h00;
            14'd279: data <= 8'h00;
            14'd280: data <= 8'h00;
            14'd281: data <= 8'h00;
            14'd282: data <= 8'h00;
            14'd283: data <= 8'h00;
            14'd284: data <= 8'h00;
            14'd285: data <= 8'h00;
            14'd286: data <= 8'h0F;
            14'd287: data <= 8'hFF;
            14'd288: data <= 8'hFF;
            14'd289: data <= 8'hFF;
            14'd290: data <= 8'hFF;
            14'd291: data <= 8'hFF;
            14'd292: data <= 8'hFF;
            14'd293: data <= 8'hFF;
            14'd294: data <= 8'hBF;
            14'd295: data <= 8'hFF;
            14'd296: data <= 8'hFF;
            14'd297: data <= 8'hFF;
            14'd298: data <= 8'hFF;
            14'd299: data <= 8'hFF;
            14'd300: data <= 8'hFF;
            14'd301: data <= 8'hFF;
            14'd302: data <= 8'hFF;
            14'd303: data <= 8'hFF;
            14'd304: data <= 8'hFF;
            14'd305: data <= 8'hFF;
            14'd306: data <= 8'hFF;
            14'd307: data <= 8'hFF;
            14'd308: data <= 8'hFF;
            14'd309: data <= 8'hFF;
            14'd310: data <= 8'hFF;
            14'd311: data <= 8'hFF;
            14'd312: data <= 8'hFF;
            14'd313: data <= 8'hF0;
            14'd314: data <= 8'h00;
            14'd315: data <= 8'h00;
            14'd316: data <= 8'h00;
            14'd317: data <= 8'h00;
            14'd318: data <= 8'h00;
            14'd319: data <= 8'h00;
            14'd320: data <= 8'h00;
            14'd321: data <= 8'h00;
            14'd322: data <= 8'h00;
            14'd323: data <= 8'h00;
            14'd324: data <= 8'h00;
            14'd325: data <= 8'h00;
            14'd326: data <= 8'h0F;
            14'd327: data <= 8'hFF;
            14'd328: data <= 8'hFF;
            14'd329: data <= 8'hFF;
            14'd330: data <= 8'hFF;
            14'd331: data <= 8'hFF;
            14'd332: data <= 8'hFF;
            14'd333: data <= 8'hFF;
            14'd334: data <= 8'hFF;
            14'd335: data <= 8'hFF;
            14'd336: data <= 8'hFF;
            14'd337: data <= 8'hFF;
            14'd338: data <= 8'hFF;
            14'd339: data <= 8'hFF;
            14'd340: data <= 8'hFF;
            14'd341: data <= 8'hFF;
            14'd342: data <= 8'hFF;
            14'd343: data <= 8'hFF;
            14'd344: data <= 8'hFF;
            14'd345: data <= 8'hFF;
            14'd346: data <= 8'hFF;
            14'd347: data <= 8'hFF;
            14'd348: data <= 8'hFF;
            14'd349: data <= 8'hFF;
            14'd350: data <= 8'hFF;
            14'd351: data <= 8'hFF;
            14'd352: data <= 8'hFF;
            14'd353: data <= 8'hF0;
            14'd354: data <= 8'h00;
            14'd355: data <= 8'h00;
            14'd356: data <= 8'h00;
            14'd357: data <= 8'h00;
            14'd358: data <= 8'h00;
            14'd359: data <= 8'h00;
            14'd360: data <= 8'h00;
            14'd361: data <= 8'h00;
            14'd362: data <= 8'h00;
            14'd363: data <= 8'h00;
            14'd364: data <= 8'h00;
            14'd365: data <= 8'h00;
            14'd366: data <= 8'h0F;
            14'd367: data <= 8'hFF;
            14'd368: data <= 8'hFF;
            14'd369: data <= 8'hFF;
            14'd370: data <= 8'hFF;
            14'd371: data <= 8'hFF;
            14'd372: data <= 8'hFF;
            14'd373: data <= 8'hFF;
            14'd374: data <= 8'hFF;
            14'd375: data <= 8'hFF;
            14'd376: data <= 8'hFF;
            14'd377: data <= 8'hFF;
            14'd378: data <= 8'hFF;
            14'd379: data <= 8'hFF;
            14'd380: data <= 8'hFF;
            14'd381: data <= 8'hFF;
            14'd382: data <= 8'hFF;
            14'd383: data <= 8'hFF;
            14'd384: data <= 8'hFF;
            14'd385: data <= 8'hFF;
            14'd386: data <= 8'hFF;
            14'd387: data <= 8'hFF;
            14'd388: data <= 8'hFF;
            14'd389: data <= 8'hFF;
            14'd390: data <= 8'hFF;
            14'd391: data <= 8'hFF;
            14'd392: data <= 8'hFF;
            14'd393: data <= 8'hF0;
            14'd394: data <= 8'h00;
            14'd395: data <= 8'h00;
            14'd396: data <= 8'h00;
            14'd397: data <= 8'h00;
            14'd398: data <= 8'h00;
            14'd399: data <= 8'h00;
            14'd400: data <= 8'h00;
            14'd401: data <= 8'h00;
            14'd402: data <= 8'h00;
            14'd403: data <= 8'h00;
            14'd404: data <= 8'h00;
            14'd405: data <= 8'h00;
            14'd406: data <= 8'h0F;
            14'd407: data <= 8'hFF;
            14'd408: data <= 8'hFF;
            14'd409: data <= 8'hFF;
            14'd410: data <= 8'hFF;
            14'd411: data <= 8'hFF;
            14'd412: data <= 8'hFF;
            14'd413: data <= 8'hFF;
            14'd414: data <= 8'hFF;
            14'd415: data <= 8'hFF;
            14'd416: data <= 8'hFF;
            14'd417: data <= 8'hFF;
            14'd418: data <= 8'hFF;
            14'd419: data <= 8'hFF;
            14'd420: data <= 8'hFF;
            14'd421: data <= 8'hFF;
            14'd422: data <= 8'hFF;
            14'd423: data <= 8'hFF;
            14'd424: data <= 8'hFF;
            14'd425: data <= 8'hFF;
            14'd426: data <= 8'hFF;
            14'd427: data <= 8'hFF;
            14'd428: data <= 8'hFF;
            14'd429: data <= 8'hFF;
            14'd430: data <= 8'hFF;
            14'd431: data <= 8'hFF;
            14'd432: data <= 8'hFF;
            14'd433: data <= 8'hF0;
            14'd434: data <= 8'h00;
            14'd435: data <= 8'h00;
            14'd436: data <= 8'h00;
            14'd437: data <= 8'h00;
            14'd438: data <= 8'h00;
            14'd439: data <= 8'h00;
            14'd440: data <= 8'h00;
            14'd441: data <= 8'h00;
            14'd442: data <= 8'h00;
            14'd443: data <= 8'h00;
            14'd444: data <= 8'h00;
            14'd445: data <= 8'h00;
            14'd446: data <= 8'h0F;
            14'd447: data <= 8'hFF;
            14'd448: data <= 8'hFF;
            14'd449: data <= 8'hFF;
            14'd450: data <= 8'hFF;
            14'd451: data <= 8'hFF;
            14'd452: data <= 8'hFF;
            14'd453: data <= 8'hFF;
            14'd454: data <= 8'hFF;
            14'd455: data <= 8'hFF;
            14'd456: data <= 8'hFF;
            14'd457: data <= 8'hFF;
            14'd458: data <= 8'hFF;
            14'd459: data <= 8'hFF;
            14'd460: data <= 8'hFF;
            14'd461: data <= 8'hFF;
            14'd462: data <= 8'h7F;
            14'd463: data <= 8'hFF;
            14'd464: data <= 8'hFF;
            14'd465: data <= 8'hFF;
            14'd466: data <= 8'hFF;
            14'd467: data <= 8'hFF;
            14'd468: data <= 8'hFF;
            14'd469: data <= 8'hFF;
            14'd470: data <= 8'hFF;
            14'd471: data <= 8'hFF;
            14'd472: data <= 8'hFF;
            14'd473: data <= 8'hF0;
            14'd474: data <= 8'h00;
            14'd475: data <= 8'h00;
            14'd476: data <= 8'h00;
            14'd477: data <= 8'h00;
            14'd478: data <= 8'h00;
            14'd479: data <= 8'h00;
            14'd480: data <= 8'h00;
            14'd481: data <= 8'h00;
            14'd482: data <= 8'h00;
            14'd483: data <= 8'h00;
            14'd484: data <= 8'h00;
            14'd485: data <= 8'h00;
            14'd486: data <= 8'h0F;
            14'd487: data <= 8'hFF;
            14'd488: data <= 8'hFF;
            14'd489: data <= 8'hFF;
            14'd490: data <= 8'hFF;
            14'd491: data <= 8'hFF;
            14'd492: data <= 8'hFF;
            14'd493: data <= 8'hFF;
            14'd494: data <= 8'hFF;
            14'd495: data <= 8'hFF;
            14'd496: data <= 8'hFF;
            14'd497: data <= 8'hFF;
            14'd498: data <= 8'hFF;
            14'd499: data <= 8'hFF;
            14'd500: data <= 8'hFF;
            14'd501: data <= 8'hFF;
            14'd502: data <= 8'hFF;
            14'd503: data <= 8'hFF;
            14'd504: data <= 8'hFF;
            14'd505: data <= 8'hFF;
            14'd506: data <= 8'hFF;
            14'd507: data <= 8'hFF;
            14'd508: data <= 8'hFF;
            14'd509: data <= 8'hFF;
            14'd510: data <= 8'hFF;
            14'd511: data <= 8'hFF;
            14'd512: data <= 8'hFF;
            14'd513: data <= 8'hF0;
            14'd514: data <= 8'h00;
            14'd515: data <= 8'h00;
            14'd516: data <= 8'h00;
            14'd517: data <= 8'h00;
            14'd518: data <= 8'h00;
            14'd519: data <= 8'h00;
            14'd520: data <= 8'h00;
            14'd521: data <= 8'h00;
            14'd522: data <= 8'h00;
            14'd523: data <= 8'h00;
            14'd524: data <= 8'h00;
            14'd525: data <= 8'h00;
            14'd526: data <= 8'h0F;
            14'd527: data <= 8'hFF;
            14'd528: data <= 8'hFF;
            14'd529: data <= 8'hFF;
            14'd530: data <= 8'hFF;
            14'd531: data <= 8'hFF;
            14'd532: data <= 8'hFF;
            14'd533: data <= 8'hFF;
            14'd534: data <= 8'hFF;
            14'd535: data <= 8'hFF;
            14'd536: data <= 8'hFF;
            14'd537: data <= 8'hFF;
            14'd538: data <= 8'hFF;
            14'd539: data <= 8'hFF;
            14'd540: data <= 8'hFF;
            14'd541: data <= 8'hFF;
            14'd542: data <= 8'hFF;
            14'd543: data <= 8'hFF;
            14'd544: data <= 8'hFF;
            14'd545: data <= 8'hFF;
            14'd546: data <= 8'hFF;
            14'd547: data <= 8'hFF;
            14'd548: data <= 8'hFF;
            14'd549: data <= 8'hFF;
            14'd550: data <= 8'hFF;
            14'd551: data <= 8'hFF;
            14'd552: data <= 8'hFF;
            14'd553: data <= 8'hF0;
            14'd554: data <= 8'h00;
            14'd555: data <= 8'h00;
            14'd556: data <= 8'h00;
            14'd557: data <= 8'h00;
            14'd558: data <= 8'h00;
            14'd559: data <= 8'h00;
            14'd560: data <= 8'h00;
            14'd561: data <= 8'h00;
            14'd562: data <= 8'h00;
            14'd563: data <= 8'h00;
            14'd564: data <= 8'h00;
            14'd565: data <= 8'h00;
            14'd566: data <= 8'h0F;
            14'd567: data <= 8'hFF;
            14'd568: data <= 8'hFF;
            14'd569: data <= 8'hFF;
            14'd570: data <= 8'hFF;
            14'd571: data <= 8'hFF;
            14'd572: data <= 8'hFF;
            14'd573: data <= 8'hFF;
            14'd574: data <= 8'hFF;
            14'd575: data <= 8'hFF;
            14'd576: data <= 8'hFF;
            14'd577: data <= 8'hFF;
            14'd578: data <= 8'hFF;
            14'd579: data <= 8'hFF;
            14'd580: data <= 8'hFF;
            14'd581: data <= 8'hFF;
            14'd582: data <= 8'hFF;
            14'd583: data <= 8'hFF;
            14'd584: data <= 8'hFF;
            14'd585: data <= 8'hFF;
            14'd586: data <= 8'hFF;
            14'd587: data <= 8'hFF;
            14'd588: data <= 8'hFF;
            14'd589: data <= 8'hFF;
            14'd590: data <= 8'hFF;
            14'd591: data <= 8'hFF;
            14'd592: data <= 8'hFF;
            14'd593: data <= 8'hF0;
            14'd594: data <= 8'h00;
            14'd595: data <= 8'h00;
            14'd596: data <= 8'h00;
            14'd597: data <= 8'h00;
            14'd598: data <= 8'h00;
            14'd599: data <= 8'h00;
            14'd600: data <= 8'h00;
            14'd601: data <= 8'h00;
            14'd602: data <= 8'h00;
            14'd603: data <= 8'h00;
            14'd604: data <= 8'h00;
            14'd605: data <= 8'h00;
            14'd606: data <= 8'h0F;
            14'd607: data <= 8'hFF;
            14'd608: data <= 8'hFF;
            14'd609: data <= 8'hFF;
            14'd610: data <= 8'hFF;
            14'd611: data <= 8'hFF;
            14'd612: data <= 8'hFF;
            14'd613: data <= 8'hFF;
            14'd614: data <= 8'hFF;
            14'd615: data <= 8'hFF;
            14'd616: data <= 8'hFF;
            14'd617: data <= 8'hFF;
            14'd618: data <= 8'hFF;
            14'd619: data <= 8'hFF;
            14'd620: data <= 8'hFF;
            14'd621: data <= 8'hFF;
            14'd622: data <= 8'hFF;
            14'd623: data <= 8'hFF;
            14'd624: data <= 8'hFF;
            14'd625: data <= 8'hFF;
            14'd626: data <= 8'hFF;
            14'd627: data <= 8'hFF;
            14'd628: data <= 8'hFF;
            14'd629: data <= 8'hFF;
            14'd630: data <= 8'hFF;
            14'd631: data <= 8'hFF;
            14'd632: data <= 8'hFF;
            14'd633: data <= 8'hF0;
            14'd634: data <= 8'h00;
            14'd635: data <= 8'h00;
            14'd636: data <= 8'h00;
            14'd637: data <= 8'h00;
            14'd638: data <= 8'h00;
            14'd639: data <= 8'h00;
            14'd640: data <= 8'h00;
            14'd641: data <= 8'h00;
            14'd642: data <= 8'h00;
            14'd643: data <= 8'h00;
            14'd644: data <= 8'h00;
            14'd645: data <= 8'h00;
            14'd646: data <= 8'h0F;
            14'd647: data <= 8'hFF;
            14'd648: data <= 8'hFF;
            14'd649: data <= 8'hFF;
            14'd650: data <= 8'hFF;
            14'd651: data <= 8'hFF;
            14'd652: data <= 8'hFF;
            14'd653: data <= 8'hFF;
            14'd654: data <= 8'hFF;
            14'd655: data <= 8'hFF;
            14'd656: data <= 8'hFF;
            14'd657: data <= 8'hFF;
            14'd658: data <= 8'hFF;
            14'd659: data <= 8'hFF;
            14'd660: data <= 8'hFF;
            14'd661: data <= 8'hFF;
            14'd662: data <= 8'hFF;
            14'd663: data <= 8'hFF;
            14'd664: data <= 8'hFF;
            14'd665: data <= 8'hFF;
            14'd666: data <= 8'hFF;
            14'd667: data <= 8'hFF;
            14'd668: data <= 8'hFF;
            14'd669: data <= 8'hFF;
            14'd670: data <= 8'hFF;
            14'd671: data <= 8'hFF;
            14'd672: data <= 8'hFF;
            14'd673: data <= 8'hF0;
            14'd674: data <= 8'h00;
            14'd675: data <= 8'h00;
            14'd676: data <= 8'h00;
            14'd677: data <= 8'h00;
            14'd678: data <= 8'h00;
            14'd679: data <= 8'h00;
            14'd680: data <= 8'h00;
            14'd681: data <= 8'h00;
            14'd682: data <= 8'h00;
            14'd683: data <= 8'h00;
            14'd684: data <= 8'h00;
            14'd685: data <= 8'h00;
            14'd686: data <= 8'h0F;
            14'd687: data <= 8'hFF;
            14'd688: data <= 8'hFF;
            14'd689: data <= 8'hFF;
            14'd690: data <= 8'hFF;
            14'd691: data <= 8'hFF;
            14'd692: data <= 8'hFF;
            14'd693: data <= 8'hFF;
            14'd694: data <= 8'hFF;
            14'd695: data <= 8'hFF;
            14'd696: data <= 8'hFF;
            14'd697: data <= 8'hFF;
            14'd698: data <= 8'hFF;
            14'd699: data <= 8'hFF;
            14'd700: data <= 8'hFF;
            14'd701: data <= 8'hFF;
            14'd702: data <= 8'hFF;
            14'd703: data <= 8'hFF;
            14'd704: data <= 8'hFF;
            14'd705: data <= 8'hFF;
            14'd706: data <= 8'hFF;
            14'd707: data <= 8'hFF;
            14'd708: data <= 8'hFF;
            14'd709: data <= 8'hFF;
            14'd710: data <= 8'hFF;
            14'd711: data <= 8'hFF;
            14'd712: data <= 8'hFF;
            14'd713: data <= 8'hF0;
            14'd714: data <= 8'h00;
            14'd715: data <= 8'h00;
            14'd716: data <= 8'h00;
            14'd717: data <= 8'h00;
            14'd718: data <= 8'h00;
            14'd719: data <= 8'h00;
            14'd720: data <= 8'h00;
            14'd721: data <= 8'h00;
            14'd722: data <= 8'h00;
            14'd723: data <= 8'h00;
            14'd724: data <= 8'h00;
            14'd725: data <= 8'h00;
            14'd726: data <= 8'h0F;
            14'd727: data <= 8'hFF;
            14'd728: data <= 8'hFF;
            14'd729: data <= 8'hFF;
            14'd730: data <= 8'hFF;
            14'd731: data <= 8'hFF;
            14'd732: data <= 8'hFF;
            14'd733: data <= 8'hFF;
            14'd734: data <= 8'hFF;
            14'd735: data <= 8'hFF;
            14'd736: data <= 8'hFF;
            14'd737: data <= 8'hFF;
            14'd738: data <= 8'hFF;
            14'd739: data <= 8'hFF;
            14'd740: data <= 8'hFF;
            14'd741: data <= 8'hFF;
            14'd742: data <= 8'hFF;
            14'd743: data <= 8'hFF;
            14'd744: data <= 8'hFF;
            14'd745: data <= 8'hFF;
            14'd746: data <= 8'hFF;
            14'd747: data <= 8'hFF;
            14'd748: data <= 8'hFF;
            14'd749: data <= 8'hFF;
            14'd750: data <= 8'hFF;
            14'd751: data <= 8'hFF;
            14'd752: data <= 8'hFF;
            14'd753: data <= 8'hF0;
            14'd754: data <= 8'h00;
            14'd755: data <= 8'h00;
            14'd756: data <= 8'h00;
            14'd757: data <= 8'h00;
            14'd758: data <= 8'h00;
            14'd759: data <= 8'h00;
            14'd760: data <= 8'h00;
            14'd761: data <= 8'h00;
            14'd762: data <= 8'h00;
            14'd763: data <= 8'h00;
            14'd764: data <= 8'h00;
            14'd765: data <= 8'h00;
            14'd766: data <= 8'h0E;
            14'd767: data <= 8'hFF;
            14'd768: data <= 8'hFF;
            14'd769: data <= 8'hFF;
            14'd770: data <= 8'hFF;
            14'd771: data <= 8'hFF;
            14'd772: data <= 8'hFF;
            14'd773: data <= 8'hFF;
            14'd774: data <= 8'hFF;
            14'd775: data <= 8'hFF;
            14'd776: data <= 8'hFF;
            14'd777: data <= 8'hFF;
            14'd778: data <= 8'hFF;
            14'd779: data <= 8'hFF;
            14'd780: data <= 8'hFF;
            14'd781: data <= 8'hFF;
            14'd782: data <= 8'hFF;
            14'd783: data <= 8'hFF;
            14'd784: data <= 8'hFF;
            14'd785: data <= 8'hFF;
            14'd786: data <= 8'hFF;
            14'd787: data <= 8'hFF;
            14'd788: data <= 8'hFF;
            14'd789: data <= 8'hFF;
            14'd790: data <= 8'hFF;
            14'd791: data <= 8'hFF;
            14'd792: data <= 8'hFF;
            14'd793: data <= 8'hF0;
            14'd794: data <= 8'h00;
            14'd795: data <= 8'h00;
            14'd796: data <= 8'h00;
            14'd797: data <= 8'h00;
            14'd798: data <= 8'h00;
            14'd799: data <= 8'h00;
            14'd800: data <= 8'h00;
            14'd801: data <= 8'h00;
            14'd802: data <= 8'h00;
            14'd803: data <= 8'h00;
            14'd804: data <= 8'h00;
            14'd805: data <= 8'h00;
            14'd806: data <= 8'h0F;
            14'd807: data <= 8'hFF;
            14'd808: data <= 8'hFF;
            14'd809: data <= 8'hFF;
            14'd810: data <= 8'hFF;
            14'd811: data <= 8'hFF;
            14'd812: data <= 8'hFF;
            14'd813: data <= 8'hFF;
            14'd814: data <= 8'hFF;
            14'd815: data <= 8'hFF;
            14'd816: data <= 8'hFF;
            14'd817: data <= 8'hBF;
            14'd818: data <= 8'hFF;
            14'd819: data <= 8'hFF;
            14'd820: data <= 8'hFF;
            14'd821: data <= 8'hFF;
            14'd822: data <= 8'hFF;
            14'd823: data <= 8'hFF;
            14'd824: data <= 8'hFF;
            14'd825: data <= 8'hFF;
            14'd826: data <= 8'hFF;
            14'd827: data <= 8'hFF;
            14'd828: data <= 8'hFF;
            14'd829: data <= 8'hFF;
            14'd830: data <= 8'hFF;
            14'd831: data <= 8'hFF;
            14'd832: data <= 8'hFF;
            14'd833: data <= 8'hF0;
            14'd834: data <= 8'h00;
            14'd835: data <= 8'h00;
            14'd836: data <= 8'h00;
            14'd837: data <= 8'h00;
            14'd838: data <= 8'h00;
            14'd839: data <= 8'h00;
            14'd840: data <= 8'h00;
            14'd841: data <= 8'h00;
            14'd842: data <= 8'h00;
            14'd843: data <= 8'h00;
            14'd844: data <= 8'h00;
            14'd845: data <= 8'h00;
            14'd846: data <= 8'h0F;
            14'd847: data <= 8'hFF;
            14'd848: data <= 8'hFF;
            14'd849: data <= 8'hFF;
            14'd850: data <= 8'hFF;
            14'd851: data <= 8'hFF;
            14'd852: data <= 8'hFF;
            14'd853: data <= 8'hFF;
            14'd854: data <= 8'hFF;
            14'd855: data <= 8'hFF;
            14'd856: data <= 8'hFF;
            14'd857: data <= 8'hFF;
            14'd858: data <= 8'hFF;
            14'd859: data <= 8'hFF;
            14'd860: data <= 8'hFF;
            14'd861: data <= 8'hFF;
            14'd862: data <= 8'hFF;
            14'd863: data <= 8'hFF;
            14'd864: data <= 8'hFF;
            14'd865: data <= 8'hFF;
            14'd866: data <= 8'hFF;
            14'd867: data <= 8'hFF;
            14'd868: data <= 8'hFF;
            14'd869: data <= 8'hFF;
            14'd870: data <= 8'hFF;
            14'd871: data <= 8'hFF;
            14'd872: data <= 8'hFF;
            14'd873: data <= 8'hF0;
            14'd874: data <= 8'h00;
            14'd875: data <= 8'h00;
            14'd876: data <= 8'h00;
            14'd877: data <= 8'h00;
            14'd878: data <= 8'h00;
            14'd879: data <= 8'h00;
            14'd880: data <= 8'h00;
            14'd881: data <= 8'h00;
            14'd882: data <= 8'h00;
            14'd883: data <= 8'h00;
            14'd884: data <= 8'h00;
            14'd885: data <= 8'h00;
            14'd886: data <= 8'h0B;
            14'd887: data <= 8'hFF;
            14'd888: data <= 8'hFF;
            14'd889: data <= 8'hFF;
            14'd890: data <= 8'hFF;
            14'd891: data <= 8'hFF;
            14'd892: data <= 8'hFF;
            14'd893: data <= 8'hFF;
            14'd894: data <= 8'hFF;
            14'd895: data <= 8'hFF;
            14'd896: data <= 8'hFF;
            14'd897: data <= 8'hFF;
            14'd898: data <= 8'hFF;
            14'd899: data <= 8'hFF;
            14'd900: data <= 8'hFF;
            14'd901: data <= 8'hFF;
            14'd902: data <= 8'hFF;
            14'd903: data <= 8'hFF;
            14'd904: data <= 8'hFF;
            14'd905: data <= 8'hFF;
            14'd906: data <= 8'hFF;
            14'd907: data <= 8'hFF;
            14'd908: data <= 8'hFF;
            14'd909: data <= 8'hFF;
            14'd910: data <= 8'hFF;
            14'd911: data <= 8'hFF;
            14'd912: data <= 8'hFF;
            14'd913: data <= 8'hF0;
            14'd914: data <= 8'h00;
            14'd915: data <= 8'h00;
            14'd916: data <= 8'h00;
            14'd917: data <= 8'h00;
            14'd918: data <= 8'h00;
            14'd919: data <= 8'h00;
            14'd920: data <= 8'h00;
            14'd921: data <= 8'h00;
            14'd922: data <= 8'h00;
            14'd923: data <= 8'h00;
            14'd924: data <= 8'h00;
            14'd925: data <= 8'h00;
            14'd926: data <= 8'h0F;
            14'd927: data <= 8'hFF;
            14'd928: data <= 8'hFF;
            14'd929: data <= 8'hFF;
            14'd930: data <= 8'hFF;
            14'd931: data <= 8'hFF;
            14'd932: data <= 8'hFF;
            14'd933: data <= 8'hFF;
            14'd934: data <= 8'hFF;
            14'd935: data <= 8'hFF;
            14'd936: data <= 8'hFF;
            14'd937: data <= 8'hFF;
            14'd938: data <= 8'hFF;
            14'd939: data <= 8'hFF;
            14'd940: data <= 8'hFF;
            14'd941: data <= 8'hFF;
            14'd942: data <= 8'hFF;
            14'd943: data <= 8'hFF;
            14'd944: data <= 8'hFF;
            14'd945: data <= 8'hFF;
            14'd946: data <= 8'hFF;
            14'd947: data <= 8'hFF;
            14'd948: data <= 8'hFF;
            14'd949: data <= 8'hFF;
            14'd950: data <= 8'hFF;
            14'd951: data <= 8'hFF;
            14'd952: data <= 8'hFF;
            14'd953: data <= 8'hF0;
            14'd954: data <= 8'h00;
            14'd955: data <= 8'h00;
            14'd956: data <= 8'h00;
            14'd957: data <= 8'h00;
            14'd958: data <= 8'h00;
            14'd959: data <= 8'h00;
            14'd960: data <= 8'h00;
            14'd961: data <= 8'h00;
            14'd962: data <= 8'h00;
            14'd963: data <= 8'h00;
            14'd964: data <= 8'h00;
            14'd965: data <= 8'h00;
            14'd966: data <= 8'h0F;
            14'd967: data <= 8'hFF;
            14'd968: data <= 8'hFF;
            14'd969: data <= 8'hFF;
            14'd970: data <= 8'hFF;
            14'd971: data <= 8'hFF;
            14'd972: data <= 8'hFF;
            14'd973: data <= 8'hFF;
            14'd974: data <= 8'hFF;
            14'd975: data <= 8'hFF;
            14'd976: data <= 8'hFF;
            14'd977: data <= 8'hFF;
            14'd978: data <= 8'hFF;
            14'd979: data <= 8'hFF;
            14'd980: data <= 8'hFF;
            14'd981: data <= 8'hFF;
            14'd982: data <= 8'hFF;
            14'd983: data <= 8'hFF;
            14'd984: data <= 8'hFF;
            14'd985: data <= 8'hFF;
            14'd986: data <= 8'hFF;
            14'd987: data <= 8'hFF;
            14'd988: data <= 8'hFF;
            14'd989: data <= 8'hFF;
            14'd990: data <= 8'hFF;
            14'd991: data <= 8'hFF;
            14'd992: data <= 8'hFF;
            14'd993: data <= 8'hF0;
            14'd994: data <= 8'h00;
            14'd995: data <= 8'h00;
            14'd996: data <= 8'h00;
            14'd997: data <= 8'h00;
            14'd998: data <= 8'h00;
            14'd999: data <= 8'h00;
            14'd1000: data <= 8'h00;
            14'd1001: data <= 8'h00;
            14'd1002: data <= 8'h00;
            14'd1003: data <= 8'h00;
            14'd1004: data <= 8'h00;
            14'd1005: data <= 8'h00;
            14'd1006: data <= 8'h0F;
            14'd1007: data <= 8'hFF;
            14'd1008: data <= 8'hFF;
            14'd1009: data <= 8'hFF;
            14'd1010: data <= 8'hFF;
            14'd1011: data <= 8'hFF;
            14'd1012: data <= 8'hFF;
            14'd1013: data <= 8'hFF;
            14'd1014: data <= 8'hFF;
            14'd1015: data <= 8'hFF;
            14'd1016: data <= 8'hFF;
            14'd1017: data <= 8'hFF;
            14'd1018: data <= 8'hFF;
            14'd1019: data <= 8'hFF;
            14'd1020: data <= 8'hFF;
            14'd1021: data <= 8'hFF;
            14'd1022: data <= 8'hFF;
            14'd1023: data <= 8'hFF;
            14'd1024: data <= 8'hFF;
            14'd1025: data <= 8'hFF;
            14'd1026: data <= 8'hFF;
            14'd1027: data <= 8'hFF;
            14'd1028: data <= 8'hFF;
            14'd1029: data <= 8'hFF;
            14'd1030: data <= 8'hFF;
            14'd1031: data <= 8'hFF;
            14'd1032: data <= 8'hFF;
            14'd1033: data <= 8'hF0;
            14'd1034: data <= 8'h00;
            14'd1035: data <= 8'h00;
            14'd1036: data <= 8'h00;
            14'd1037: data <= 8'h00;
            14'd1038: data <= 8'h00;
            14'd1039: data <= 8'h00;
            14'd1040: data <= 8'h00;
            14'd1041: data <= 8'h00;
            14'd1042: data <= 8'h00;
            14'd1043: data <= 8'h00;
            14'd1044: data <= 8'h00;
            14'd1045: data <= 8'h00;
            14'd1046: data <= 8'h0F;
            14'd1047: data <= 8'hFF;
            14'd1048: data <= 8'hFF;
            14'd1049: data <= 8'hFF;
            14'd1050: data <= 8'hFF;
            14'd1051: data <= 8'hFF;
            14'd1052: data <= 8'hFF;
            14'd1053: data <= 8'hFF;
            14'd1054: data <= 8'hFF;
            14'd1055: data <= 8'hFF;
            14'd1056: data <= 8'hFF;
            14'd1057: data <= 8'hFF;
            14'd1058: data <= 8'hFF;
            14'd1059: data <= 8'hFF;
            14'd1060: data <= 8'hFF;
            14'd1061: data <= 8'hFF;
            14'd1062: data <= 8'hFF;
            14'd1063: data <= 8'hFF;
            14'd1064: data <= 8'hFF;
            14'd1065: data <= 8'hFF;
            14'd1066: data <= 8'hFF;
            14'd1067: data <= 8'hFF;
            14'd1068: data <= 8'hFF;
            14'd1069: data <= 8'hFF;
            14'd1070: data <= 8'hFF;
            14'd1071: data <= 8'hFF;
            14'd1072: data <= 8'hFF;
            14'd1073: data <= 8'hF0;
            14'd1074: data <= 8'h00;
            14'd1075: data <= 8'h00;
            14'd1076: data <= 8'h00;
            14'd1077: data <= 8'h00;
            14'd1078: data <= 8'h00;
            14'd1079: data <= 8'h00;
            14'd1080: data <= 8'h00;
            14'd1081: data <= 8'h00;
            14'd1082: data <= 8'h00;
            14'd1083: data <= 8'h00;
            14'd1084: data <= 8'h00;
            14'd1085: data <= 8'h00;
            14'd1086: data <= 8'h0F;
            14'd1087: data <= 8'hFF;
            14'd1088: data <= 8'hFF;
            14'd1089: data <= 8'hFF;
            14'd1090: data <= 8'hFF;
            14'd1091: data <= 8'hFF;
            14'd1092: data <= 8'hFF;
            14'd1093: data <= 8'hFF;
            14'd1094: data <= 8'hFF;
            14'd1095: data <= 8'hFF;
            14'd1096: data <= 8'hFF;
            14'd1097: data <= 8'hFF;
            14'd1098: data <= 8'hFF;
            14'd1099: data <= 8'hFF;
            14'd1100: data <= 8'hFF;
            14'd1101: data <= 8'hFF;
            14'd1102: data <= 8'hFF;
            14'd1103: data <= 8'hFF;
            14'd1104: data <= 8'hFF;
            14'd1105: data <= 8'hFF;
            14'd1106: data <= 8'hFF;
            14'd1107: data <= 8'hFF;
            14'd1108: data <= 8'hFF;
            14'd1109: data <= 8'hFF;
            14'd1110: data <= 8'hFF;
            14'd1111: data <= 8'hFF;
            14'd1112: data <= 8'hFF;
            14'd1113: data <= 8'hF0;
            14'd1114: data <= 8'h00;
            14'd1115: data <= 8'h00;
            14'd1116: data <= 8'h00;
            14'd1117: data <= 8'h00;
            14'd1118: data <= 8'h00;
            14'd1119: data <= 8'h00;
            14'd1120: data <= 8'h00;
            14'd1121: data <= 8'h00;
            14'd1122: data <= 8'h00;
            14'd1123: data <= 8'h00;
            14'd1124: data <= 8'h00;
            14'd1125: data <= 8'h00;
            14'd1126: data <= 8'h0F;
            14'd1127: data <= 8'hFF;
            14'd1128: data <= 8'hFF;
            14'd1129: data <= 8'hFF;
            14'd1130: data <= 8'hFF;
            14'd1131: data <= 8'hFF;
            14'd1132: data <= 8'hFF;
            14'd1133: data <= 8'hFF;
            14'd1134: data <= 8'hFF;
            14'd1135: data <= 8'hFF;
            14'd1136: data <= 8'hFF;
            14'd1137: data <= 8'hFF;
            14'd1138: data <= 8'hFF;
            14'd1139: data <= 8'hFF;
            14'd1140: data <= 8'hFF;
            14'd1141: data <= 8'hFF;
            14'd1142: data <= 8'hFF;
            14'd1143: data <= 8'hFF;
            14'd1144: data <= 8'hFF;
            14'd1145: data <= 8'hFF;
            14'd1146: data <= 8'hFF;
            14'd1147: data <= 8'hFF;
            14'd1148: data <= 8'hFF;
            14'd1149: data <= 8'hFF;
            14'd1150: data <= 8'hFF;
            14'd1151: data <= 8'hFF;
            14'd1152: data <= 8'hFF;
            14'd1153: data <= 8'hF0;
            14'd1154: data <= 8'h00;
            14'd1155: data <= 8'h00;
            14'd1156: data <= 8'h00;
            14'd1157: data <= 8'h00;
            14'd1158: data <= 8'h00;
            14'd1159: data <= 8'h00;
            14'd1160: data <= 8'h00;
            14'd1161: data <= 8'h00;
            14'd1162: data <= 8'h00;
            14'd1163: data <= 8'h00;
            14'd1164: data <= 8'h00;
            14'd1165: data <= 8'h00;
            14'd1166: data <= 8'h0F;
            14'd1167: data <= 8'hFF;
            14'd1168: data <= 8'hFF;
            14'd1169: data <= 8'hFF;
            14'd1170: data <= 8'hFF;
            14'd1171: data <= 8'hFF;
            14'd1172: data <= 8'hFF;
            14'd1173: data <= 8'hFF;
            14'd1174: data <= 8'hFF;
            14'd1175: data <= 8'hFF;
            14'd1176: data <= 8'hFF;
            14'd1177: data <= 8'hFF;
            14'd1178: data <= 8'hFF;
            14'd1179: data <= 8'hFF;
            14'd1180: data <= 8'hFF;
            14'd1181: data <= 8'hFF;
            14'd1182: data <= 8'hFF;
            14'd1183: data <= 8'hFF;
            14'd1184: data <= 8'hFF;
            14'd1185: data <= 8'hFF;
            14'd1186: data <= 8'hFF;
            14'd1187: data <= 8'hFF;
            14'd1188: data <= 8'hFF;
            14'd1189: data <= 8'hFF;
            14'd1190: data <= 8'hFF;
            14'd1191: data <= 8'hFF;
            14'd1192: data <= 8'hFF;
            14'd1193: data <= 8'hF0;
            14'd1194: data <= 8'h00;
            14'd1195: data <= 8'h00;
            14'd1196: data <= 8'h00;
            14'd1197: data <= 8'h00;
            14'd1198: data <= 8'h00;
            14'd1199: data <= 8'h00;
            14'd1200: data <= 8'h00;
            14'd1201: data <= 8'h00;
            14'd1202: data <= 8'h00;
            14'd1203: data <= 8'h00;
            14'd1204: data <= 8'h00;
            14'd1205: data <= 8'h00;
            14'd1206: data <= 8'h0F;
            14'd1207: data <= 8'hFF;
            14'd1208: data <= 8'hFF;
            14'd1209: data <= 8'hFF;
            14'd1210: data <= 8'hFF;
            14'd1211: data <= 8'hFF;
            14'd1212: data <= 8'hFF;
            14'd1213: data <= 8'hFF;
            14'd1214: data <= 8'hFF;
            14'd1215: data <= 8'hFF;
            14'd1216: data <= 8'hFF;
            14'd1217: data <= 8'hFF;
            14'd1218: data <= 8'hFF;
            14'd1219: data <= 8'hFF;
            14'd1220: data <= 8'hEF;
            14'd1221: data <= 8'hFF;
            14'd1222: data <= 8'hFF;
            14'd1223: data <= 8'hFF;
            14'd1224: data <= 8'hFF;
            14'd1225: data <= 8'hFF;
            14'd1226: data <= 8'hFF;
            14'd1227: data <= 8'hFF;
            14'd1228: data <= 8'hFF;
            14'd1229: data <= 8'hFF;
            14'd1230: data <= 8'hFF;
            14'd1231: data <= 8'hFF;
            14'd1232: data <= 8'hFF;
            14'd1233: data <= 8'hF0;
            14'd1234: data <= 8'h00;
            14'd1235: data <= 8'h00;
            14'd1236: data <= 8'h00;
            14'd1237: data <= 8'h00;
            14'd1238: data <= 8'h00;
            14'd1239: data <= 8'h00;
            14'd1240: data <= 8'h00;
            14'd1241: data <= 8'h00;
            14'd1242: data <= 8'h00;
            14'd1243: data <= 8'h00;
            14'd1244: data <= 8'h00;
            14'd1245: data <= 8'h00;
            14'd1246: data <= 8'h0F;
            14'd1247: data <= 8'hFF;
            14'd1248: data <= 8'hFF;
            14'd1249: data <= 8'hFF;
            14'd1250: data <= 8'hFF;
            14'd1251: data <= 8'hFF;
            14'd1252: data <= 8'hFF;
            14'd1253: data <= 8'hFF;
            14'd1254: data <= 8'hFF;
            14'd1255: data <= 8'hFF;
            14'd1256: data <= 8'hFF;
            14'd1257: data <= 8'hFF;
            14'd1258: data <= 8'hFF;
            14'd1259: data <= 8'hFF;
            14'd1260: data <= 8'hFF;
            14'd1261: data <= 8'hFF;
            14'd1262: data <= 8'hFF;
            14'd1263: data <= 8'hFF;
            14'd1264: data <= 8'hFF;
            14'd1265: data <= 8'hFF;
            14'd1266: data <= 8'hFF;
            14'd1267: data <= 8'hFF;
            14'd1268: data <= 8'hFF;
            14'd1269: data <= 8'hFF;
            14'd1270: data <= 8'hFF;
            14'd1271: data <= 8'hFF;
            14'd1272: data <= 8'hFF;
            14'd1273: data <= 8'hF0;
            14'd1274: data <= 8'h00;
            14'd1275: data <= 8'h00;
            14'd1276: data <= 8'h00;
            14'd1277: data <= 8'h00;
            14'd1278: data <= 8'h00;
            14'd1279: data <= 8'h00;
            14'd1280: data <= 8'h00;
            14'd1281: data <= 8'h00;
            14'd1282: data <= 8'h00;
            14'd1283: data <= 8'h00;
            14'd1284: data <= 8'h00;
            14'd1285: data <= 8'h00;
            14'd1286: data <= 8'h0F;
            14'd1287: data <= 8'hFF;
            14'd1288: data <= 8'hFF;
            14'd1289: data <= 8'hFF;
            14'd1290: data <= 8'hFF;
            14'd1291: data <= 8'hFF;
            14'd1292: data <= 8'hFF;
            14'd1293: data <= 8'hFF;
            14'd1294: data <= 8'hFF;
            14'd1295: data <= 8'hFF;
            14'd1296: data <= 8'hFF;
            14'd1297: data <= 8'hFF;
            14'd1298: data <= 8'hFF;
            14'd1299: data <= 8'hFF;
            14'd1300: data <= 8'hFF;
            14'd1301: data <= 8'hFF;
            14'd1302: data <= 8'hFF;
            14'd1303: data <= 8'hFF;
            14'd1304: data <= 8'hFF;
            14'd1305: data <= 8'hFF;
            14'd1306: data <= 8'hFF;
            14'd1307: data <= 8'hFF;
            14'd1308: data <= 8'hFF;
            14'd1309: data <= 8'hFF;
            14'd1310: data <= 8'hFF;
            14'd1311: data <= 8'hFF;
            14'd1312: data <= 8'hFF;
            14'd1313: data <= 8'hF0;
            14'd1314: data <= 8'h00;
            14'd1315: data <= 8'h00;
            14'd1316: data <= 8'h00;
            14'd1317: data <= 8'h00;
            14'd1318: data <= 8'h00;
            14'd1319: data <= 8'h00;
            14'd1320: data <= 8'h00;
            14'd1321: data <= 8'h00;
            14'd1322: data <= 8'h00;
            14'd1323: data <= 8'h00;
            14'd1324: data <= 8'h00;
            14'd1325: data <= 8'h00;
            14'd1326: data <= 8'h0F;
            14'd1327: data <= 8'hFF;
            14'd1328: data <= 8'hFF;
            14'd1329: data <= 8'hFF;
            14'd1330: data <= 8'hFF;
            14'd1331: data <= 8'hFF;
            14'd1332: data <= 8'hFF;
            14'd1333: data <= 8'hFF;
            14'd1334: data <= 8'hFF;
            14'd1335: data <= 8'hFF;
            14'd1336: data <= 8'hFF;
            14'd1337: data <= 8'hFF;
            14'd1338: data <= 8'hFF;
            14'd1339: data <= 8'hFF;
            14'd1340: data <= 8'hFF;
            14'd1341: data <= 8'hFF;
            14'd1342: data <= 8'hFF;
            14'd1343: data <= 8'hFF;
            14'd1344: data <= 8'hFF;
            14'd1345: data <= 8'hFF;
            14'd1346: data <= 8'hFF;
            14'd1347: data <= 8'hFF;
            14'd1348: data <= 8'hFF;
            14'd1349: data <= 8'hFF;
            14'd1350: data <= 8'hFF;
            14'd1351: data <= 8'hFF;
            14'd1352: data <= 8'hFF;
            14'd1353: data <= 8'hF0;
            14'd1354: data <= 8'h00;
            14'd1355: data <= 8'h00;
            14'd1356: data <= 8'h00;
            14'd1357: data <= 8'h00;
            14'd1358: data <= 8'h00;
            14'd1359: data <= 8'h00;
            14'd1360: data <= 8'h00;
            14'd1361: data <= 8'h00;
            14'd1362: data <= 8'h00;
            14'd1363: data <= 8'h00;
            14'd1364: data <= 8'h00;
            14'd1365: data <= 8'h00;
            14'd1366: data <= 8'h0F;
            14'd1367: data <= 8'hFF;
            14'd1368: data <= 8'hFF;
            14'd1369: data <= 8'hFF;
            14'd1370: data <= 8'hFF;
            14'd1371: data <= 8'hFF;
            14'd1372: data <= 8'hFF;
            14'd1373: data <= 8'hFF;
            14'd1374: data <= 8'hFF;
            14'd1375: data <= 8'hFF;
            14'd1376: data <= 8'hFF;
            14'd1377: data <= 8'hFF;
            14'd1378: data <= 8'hFF;
            14'd1379: data <= 8'hFF;
            14'd1380: data <= 8'hFF;
            14'd1381: data <= 8'hFF;
            14'd1382: data <= 8'hFF;
            14'd1383: data <= 8'hFF;
            14'd1384: data <= 8'hFF;
            14'd1385: data <= 8'hFF;
            14'd1386: data <= 8'hFF;
            14'd1387: data <= 8'hFF;
            14'd1388: data <= 8'hFF;
            14'd1389: data <= 8'hFF;
            14'd1390: data <= 8'hFF;
            14'd1391: data <= 8'hFF;
            14'd1392: data <= 8'hFF;
            14'd1393: data <= 8'hF0;
            14'd1394: data <= 8'h00;
            14'd1395: data <= 8'h00;
            14'd1396: data <= 8'h00;
            14'd1397: data <= 8'h00;
            14'd1398: data <= 8'h00;
            14'd1399: data <= 8'h00;
            14'd1400: data <= 8'h00;
            14'd1401: data <= 8'h00;
            14'd1402: data <= 8'h00;
            14'd1403: data <= 8'h00;
            14'd1404: data <= 8'h00;
            14'd1405: data <= 8'h00;
            14'd1406: data <= 8'h0F;
            14'd1407: data <= 8'hFF;
            14'd1408: data <= 8'hFF;
            14'd1409: data <= 8'hFF;
            14'd1410: data <= 8'hFF;
            14'd1411: data <= 8'hFF;
            14'd1412: data <= 8'hFF;
            14'd1413: data <= 8'hFF;
            14'd1414: data <= 8'hFF;
            14'd1415: data <= 8'hFF;
            14'd1416: data <= 8'hFF;
            14'd1417: data <= 8'hFF;
            14'd1418: data <= 8'hFF;
            14'd1419: data <= 8'hFF;
            14'd1420: data <= 8'hFF;
            14'd1421: data <= 8'hFF;
            14'd1422: data <= 8'hFF;
            14'd1423: data <= 8'hFF;
            14'd1424: data <= 8'hFF;
            14'd1425: data <= 8'hFF;
            14'd1426: data <= 8'hFF;
            14'd1427: data <= 8'hFF;
            14'd1428: data <= 8'hFF;
            14'd1429: data <= 8'hFF;
            14'd1430: data <= 8'hFF;
            14'd1431: data <= 8'hFF;
            14'd1432: data <= 8'hFF;
            14'd1433: data <= 8'hF0;
            14'd1434: data <= 8'h00;
            14'd1435: data <= 8'h00;
            14'd1436: data <= 8'h00;
            14'd1437: data <= 8'h00;
            14'd1438: data <= 8'h00;
            14'd1439: data <= 8'h00;
            14'd1440: data <= 8'h00;
            14'd1441: data <= 8'h00;
            14'd1442: data <= 8'h00;
            14'd1443: data <= 8'h00;
            14'd1444: data <= 8'h00;
            14'd1445: data <= 8'h00;
            14'd1446: data <= 8'h0F;
            14'd1447: data <= 8'hFF;
            14'd1448: data <= 8'hFF;
            14'd1449: data <= 8'hFF;
            14'd1450: data <= 8'hFF;
            14'd1451: data <= 8'hFF;
            14'd1452: data <= 8'hFF;
            14'd1453: data <= 8'hFF;
            14'd1454: data <= 8'hFF;
            14'd1455: data <= 8'hFF;
            14'd1456: data <= 8'hFF;
            14'd1457: data <= 8'hFF;
            14'd1458: data <= 8'hFF;
            14'd1459: data <= 8'hFF;
            14'd1460: data <= 8'hFF;
            14'd1461: data <= 8'hFF;
            14'd1462: data <= 8'hFF;
            14'd1463: data <= 8'hFF;
            14'd1464: data <= 8'hFF;
            14'd1465: data <= 8'hFF;
            14'd1466: data <= 8'hFF;
            14'd1467: data <= 8'hFF;
            14'd1468: data <= 8'hFF;
            14'd1469: data <= 8'hFF;
            14'd1470: data <= 8'hFF;
            14'd1471: data <= 8'hFF;
            14'd1472: data <= 8'hFF;
            14'd1473: data <= 8'hF0;
            14'd1474: data <= 8'h00;
            14'd1475: data <= 8'h00;
            14'd1476: data <= 8'h00;
            14'd1477: data <= 8'h00;
            14'd1478: data <= 8'h00;
            14'd1479: data <= 8'h00;
            14'd1480: data <= 8'h00;
            14'd1481: data <= 8'h00;
            14'd1482: data <= 8'h00;
            14'd1483: data <= 8'h00;
            14'd1484: data <= 8'h00;
            14'd1485: data <= 8'h00;
            14'd1486: data <= 8'h0F;
            14'd1487: data <= 8'hFF;
            14'd1488: data <= 8'hFF;
            14'd1489: data <= 8'hFF;
            14'd1490: data <= 8'hFF;
            14'd1491: data <= 8'hFF;
            14'd1492: data <= 8'hFF;
            14'd1493: data <= 8'hFF;
            14'd1494: data <= 8'hFF;
            14'd1495: data <= 8'hFF;
            14'd1496: data <= 8'hFF;
            14'd1497: data <= 8'hFF;
            14'd1498: data <= 8'hFF;
            14'd1499: data <= 8'hFF;
            14'd1500: data <= 8'hFF;
            14'd1501: data <= 8'hFF;
            14'd1502: data <= 8'hFF;
            14'd1503: data <= 8'hFF;
            14'd1504: data <= 8'hFF;
            14'd1505: data <= 8'hFF;
            14'd1506: data <= 8'hFF;
            14'd1507: data <= 8'hFF;
            14'd1508: data <= 8'hFF;
            14'd1509: data <= 8'hFF;
            14'd1510: data <= 8'hFF;
            14'd1511: data <= 8'hFF;
            14'd1512: data <= 8'hFF;
            14'd1513: data <= 8'hF0;
            14'd1514: data <= 8'h00;
            14'd1515: data <= 8'h00;
            14'd1516: data <= 8'h00;
            14'd1517: data <= 8'h00;
            14'd1518: data <= 8'h00;
            14'd1519: data <= 8'h00;
            14'd1520: data <= 8'h00;
            14'd1521: data <= 8'h00;
            14'd1522: data <= 8'h00;
            14'd1523: data <= 8'h00;
            14'd1524: data <= 8'h00;
            14'd1525: data <= 8'h00;
            14'd1526: data <= 8'h0F;
            14'd1527: data <= 8'hFF;
            14'd1528: data <= 8'hFF;
            14'd1529: data <= 8'hFF;
            14'd1530: data <= 8'h7F;
            14'd1531: data <= 8'hFF;
            14'd1532: data <= 8'hFF;
            14'd1533: data <= 8'hFF;
            14'd1534: data <= 8'hFF;
            14'd1535: data <= 8'hFF;
            14'd1536: data <= 8'hFF;
            14'd1537: data <= 8'hFF;
            14'd1538: data <= 8'hFF;
            14'd1539: data <= 8'hFF;
            14'd1540: data <= 8'hFF;
            14'd1541: data <= 8'hFF;
            14'd1542: data <= 8'hFF;
            14'd1543: data <= 8'hFF;
            14'd1544: data <= 8'hFF;
            14'd1545: data <= 8'hFF;
            14'd1546: data <= 8'hFF;
            14'd1547: data <= 8'hFF;
            14'd1548: data <= 8'hFF;
            14'd1549: data <= 8'hFF;
            14'd1550: data <= 8'hFF;
            14'd1551: data <= 8'hFF;
            14'd1552: data <= 8'hFF;
            14'd1553: data <= 8'hF0;
            14'd1554: data <= 8'h00;
            14'd1555: data <= 8'h00;
            14'd1556: data <= 8'h00;
            14'd1557: data <= 8'h00;
            14'd1558: data <= 8'h00;
            14'd1559: data <= 8'h00;
            14'd1560: data <= 8'h00;
            14'd1561: data <= 8'h00;
            14'd1562: data <= 8'h00;
            14'd1563: data <= 8'h00;
            14'd1564: data <= 8'h00;
            14'd1565: data <= 8'h00;
            14'd1566: data <= 8'h0F;
            14'd1567: data <= 8'hFF;
            14'd1568: data <= 8'hFF;
            14'd1569: data <= 8'hFF;
            14'd1570: data <= 8'hFF;
            14'd1571: data <= 8'hFF;
            14'd1572: data <= 8'hFF;
            14'd1573: data <= 8'hFF;
            14'd1574: data <= 8'hFF;
            14'd1575: data <= 8'hFF;
            14'd1576: data <= 8'hFF;
            14'd1577: data <= 8'hFF;
            14'd1578: data <= 8'hFF;
            14'd1579: data <= 8'hFF;
            14'd1580: data <= 8'hFF;
            14'd1581: data <= 8'hFF;
            14'd1582: data <= 8'hFF;
            14'd1583: data <= 8'hFF;
            14'd1584: data <= 8'hFF;
            14'd1585: data <= 8'hFF;
            14'd1586: data <= 8'hFF;
            14'd1587: data <= 8'hFF;
            14'd1588: data <= 8'hFF;
            14'd1589: data <= 8'hFF;
            14'd1590: data <= 8'hFF;
            14'd1591: data <= 8'hFF;
            14'd1592: data <= 8'hFF;
            14'd1593: data <= 8'hF0;
            14'd1594: data <= 8'h00;
            14'd1595: data <= 8'h00;
            14'd1596: data <= 8'h00;
            14'd1597: data <= 8'h00;
            14'd1598: data <= 8'h00;
            14'd1599: data <= 8'h00;
            14'd1600: data <= 8'h00;
            14'd1601: data <= 8'h00;
            14'd1602: data <= 8'h00;
            14'd1603: data <= 8'h00;
            14'd1604: data <= 8'h00;
            14'd1605: data <= 8'h00;
            14'd1606: data <= 8'h0F;
            14'd1607: data <= 8'hFF;
            14'd1608: data <= 8'hFF;
            14'd1609: data <= 8'hFF;
            14'd1610: data <= 8'hFF;
            14'd1611: data <= 8'hFF;
            14'd1612: data <= 8'hFF;
            14'd1613: data <= 8'hFF;
            14'd1614: data <= 8'hFF;
            14'd1615: data <= 8'hFF;
            14'd1616: data <= 8'hFF;
            14'd1617: data <= 8'hFF;
            14'd1618: data <= 8'hFF;
            14'd1619: data <= 8'hFF;
            14'd1620: data <= 8'hFF;
            14'd1621: data <= 8'hFF;
            14'd1622: data <= 8'hFF;
            14'd1623: data <= 8'hFF;
            14'd1624: data <= 8'hFF;
            14'd1625: data <= 8'hFF;
            14'd1626: data <= 8'hFF;
            14'd1627: data <= 8'hFF;
            14'd1628: data <= 8'hFF;
            14'd1629: data <= 8'hFF;
            14'd1630: data <= 8'hFF;
            14'd1631: data <= 8'hFF;
            14'd1632: data <= 8'hFF;
            14'd1633: data <= 8'hF0;
            14'd1634: data <= 8'h00;
            14'd1635: data <= 8'h00;
            14'd1636: data <= 8'h00;
            14'd1637: data <= 8'h00;
            14'd1638: data <= 8'h00;
            14'd1639: data <= 8'h00;
            14'd1640: data <= 8'h00;
            14'd1641: data <= 8'h00;
            14'd1642: data <= 8'h00;
            14'd1643: data <= 8'h00;
            14'd1644: data <= 8'h00;
            14'd1645: data <= 8'h00;
            14'd1646: data <= 8'h0F;
            14'd1647: data <= 8'hFF;
            14'd1648: data <= 8'hFF;
            14'd1649: data <= 8'hFF;
            14'd1650: data <= 8'hFF;
            14'd1651: data <= 8'hFF;
            14'd1652: data <= 8'hFF;
            14'd1653: data <= 8'hFF;
            14'd1654: data <= 8'hFF;
            14'd1655: data <= 8'hFF;
            14'd1656: data <= 8'hFF;
            14'd1657: data <= 8'hFF;
            14'd1658: data <= 8'hFF;
            14'd1659: data <= 8'hFF;
            14'd1660: data <= 8'hFF;
            14'd1661: data <= 8'hFF;
            14'd1662: data <= 8'hFF;
            14'd1663: data <= 8'hFF;
            14'd1664: data <= 8'hFF;
            14'd1665: data <= 8'hFF;
            14'd1666: data <= 8'hFF;
            14'd1667: data <= 8'hFF;
            14'd1668: data <= 8'hFF;
            14'd1669: data <= 8'hFF;
            14'd1670: data <= 8'hFF;
            14'd1671: data <= 8'hFF;
            14'd1672: data <= 8'hFF;
            14'd1673: data <= 8'hF0;
            14'd1674: data <= 8'h00;
            14'd1675: data <= 8'h00;
            14'd1676: data <= 8'h00;
            14'd1677: data <= 8'h00;
            14'd1678: data <= 8'h00;
            14'd1679: data <= 8'h00;
            14'd1680: data <= 8'h00;
            14'd1681: data <= 8'h00;
            14'd1682: data <= 8'h00;
            14'd1683: data <= 8'h00;
            14'd1684: data <= 8'h00;
            14'd1685: data <= 8'h00;
            14'd1686: data <= 8'h0F;
            14'd1687: data <= 8'hFF;
            14'd1688: data <= 8'hFF;
            14'd1689: data <= 8'hFF;
            14'd1690: data <= 8'hFF;
            14'd1691: data <= 8'hFF;
            14'd1692: data <= 8'hFF;
            14'd1693: data <= 8'hFF;
            14'd1694: data <= 8'hFF;
            14'd1695: data <= 8'hFF;
            14'd1696: data <= 8'hFF;
            14'd1697: data <= 8'hFF;
            14'd1698: data <= 8'hFF;
            14'd1699: data <= 8'hFF;
            14'd1700: data <= 8'hFF;
            14'd1701: data <= 8'hFF;
            14'd1702: data <= 8'hFF;
            14'd1703: data <= 8'hFF;
            14'd1704: data <= 8'hFF;
            14'd1705: data <= 8'hFF;
            14'd1706: data <= 8'hFF;
            14'd1707: data <= 8'hFF;
            14'd1708: data <= 8'hFF;
            14'd1709: data <= 8'hFF;
            14'd1710: data <= 8'hFF;
            14'd1711: data <= 8'hFF;
            14'd1712: data <= 8'hFF;
            14'd1713: data <= 8'hF0;
            14'd1714: data <= 8'h00;
            14'd1715: data <= 8'h00;
            14'd1716: data <= 8'h00;
            14'd1717: data <= 8'h00;
            14'd1718: data <= 8'h00;
            14'd1719: data <= 8'h00;
            14'd1720: data <= 8'h00;
            14'd1721: data <= 8'h00;
            14'd1722: data <= 8'h00;
            14'd1723: data <= 8'h00;
            14'd1724: data <= 8'h00;
            14'd1725: data <= 8'h00;
            14'd1726: data <= 8'h0F;
            14'd1727: data <= 8'hFF;
            14'd1728: data <= 8'hFF;
            14'd1729: data <= 8'hFF;
            14'd1730: data <= 8'hFF;
            14'd1731: data <= 8'hFF;
            14'd1732: data <= 8'hFF;
            14'd1733: data <= 8'hFF;
            14'd1734: data <= 8'hFF;
            14'd1735: data <= 8'hFF;
            14'd1736: data <= 8'hFF;
            14'd1737: data <= 8'hFF;
            14'd1738: data <= 8'hFF;
            14'd1739: data <= 8'hFF;
            14'd1740: data <= 8'hFF;
            14'd1741: data <= 8'hFF;
            14'd1742: data <= 8'hFF;
            14'd1743: data <= 8'hFF;
            14'd1744: data <= 8'hFF;
            14'd1745: data <= 8'hFF;
            14'd1746: data <= 8'hFF;
            14'd1747: data <= 8'hFF;
            14'd1748: data <= 8'hFF;
            14'd1749: data <= 8'hFF;
            14'd1750: data <= 8'hFF;
            14'd1751: data <= 8'hFF;
            14'd1752: data <= 8'hFF;
            14'd1753: data <= 8'hF0;
            14'd1754: data <= 8'h00;
            14'd1755: data <= 8'h00;
            14'd1756: data <= 8'h00;
            14'd1757: data <= 8'h00;
            14'd1758: data <= 8'h00;
            14'd1759: data <= 8'h00;
            14'd1760: data <= 8'h00;
            14'd1761: data <= 8'h00;
            14'd1762: data <= 8'h00;
            14'd1763: data <= 8'h00;
            14'd1764: data <= 8'h00;
            14'd1765: data <= 8'h00;
            14'd1766: data <= 8'h0F;
            14'd1767: data <= 8'hFF;
            14'd1768: data <= 8'hFF;
            14'd1769: data <= 8'hFF;
            14'd1770: data <= 8'hFF;
            14'd1771: data <= 8'hFF;
            14'd1772: data <= 8'hFF;
            14'd1773: data <= 8'hFF;
            14'd1774: data <= 8'hFF;
            14'd1775: data <= 8'hFF;
            14'd1776: data <= 8'hFF;
            14'd1777: data <= 8'hFF;
            14'd1778: data <= 8'hFF;
            14'd1779: data <= 8'hFF;
            14'd1780: data <= 8'hFF;
            14'd1781: data <= 8'hFF;
            14'd1782: data <= 8'hFF;
            14'd1783: data <= 8'hFF;
            14'd1784: data <= 8'hFF;
            14'd1785: data <= 8'hFF;
            14'd1786: data <= 8'hFF;
            14'd1787: data <= 8'hFF;
            14'd1788: data <= 8'hFF;
            14'd1789: data <= 8'hFF;
            14'd1790: data <= 8'hFF;
            14'd1791: data <= 8'hFF;
            14'd1792: data <= 8'hFF;
            14'd1793: data <= 8'hF0;
            14'd1794: data <= 8'h00;
            14'd1795: data <= 8'h00;
            14'd1796: data <= 8'h00;
            14'd1797: data <= 8'h00;
            14'd1798: data <= 8'h00;
            14'd1799: data <= 8'h00;
            14'd1800: data <= 8'h00;
            14'd1801: data <= 8'h00;
            14'd1802: data <= 8'h00;
            14'd1803: data <= 8'h00;
            14'd1804: data <= 8'h00;
            14'd1805: data <= 8'h00;
            14'd1806: data <= 8'h0F;
            14'd1807: data <= 8'hFF;
            14'd1808: data <= 8'hFF;
            14'd1809: data <= 8'hFF;
            14'd1810: data <= 8'hFF;
            14'd1811: data <= 8'hFF;
            14'd1812: data <= 8'hFF;
            14'd1813: data <= 8'hFF;
            14'd1814: data <= 8'hFF;
            14'd1815: data <= 8'hFF;
            14'd1816: data <= 8'hFF;
            14'd1817: data <= 8'hFF;
            14'd1818: data <= 8'hFF;
            14'd1819: data <= 8'hFF;
            14'd1820: data <= 8'hFF;
            14'd1821: data <= 8'hFF;
            14'd1822: data <= 8'hFF;
            14'd1823: data <= 8'hFF;
            14'd1824: data <= 8'hFF;
            14'd1825: data <= 8'hFF;
            14'd1826: data <= 8'hFF;
            14'd1827: data <= 8'hFF;
            14'd1828: data <= 8'hFF;
            14'd1829: data <= 8'hFF;
            14'd1830: data <= 8'hFF;
            14'd1831: data <= 8'hFF;
            14'd1832: data <= 8'hFF;
            14'd1833: data <= 8'hF0;
            14'd1834: data <= 8'h00;
            14'd1835: data <= 8'h00;
            14'd1836: data <= 8'h00;
            14'd1837: data <= 8'h00;
            14'd1838: data <= 8'h00;
            14'd1839: data <= 8'h00;
            14'd1840: data <= 8'h00;
            14'd1841: data <= 8'h00;
            14'd1842: data <= 8'h00;
            14'd1843: data <= 8'h00;
            14'd1844: data <= 8'h00;
            14'd1845: data <= 8'h00;
            14'd1846: data <= 8'h0F;
            14'd1847: data <= 8'hFF;
            14'd1848: data <= 8'hFF;
            14'd1849: data <= 8'hFF;
            14'd1850: data <= 8'hFF;
            14'd1851: data <= 8'hFF;
            14'd1852: data <= 8'hFF;
            14'd1853: data <= 8'hFF;
            14'd1854: data <= 8'hFF;
            14'd1855: data <= 8'hFF;
            14'd1856: data <= 8'hFF;
            14'd1857: data <= 8'hFF;
            14'd1858: data <= 8'hFF;
            14'd1859: data <= 8'hFF;
            14'd1860: data <= 8'hFF;
            14'd1861: data <= 8'hFF;
            14'd1862: data <= 8'hFF;
            14'd1863: data <= 8'hFF;
            14'd1864: data <= 8'hFF;
            14'd1865: data <= 8'hFF;
            14'd1866: data <= 8'hFF;
            14'd1867: data <= 8'hFF;
            14'd1868: data <= 8'hFF;
            14'd1869: data <= 8'hFF;
            14'd1870: data <= 8'hFF;
            14'd1871: data <= 8'hFF;
            14'd1872: data <= 8'hFF;
            14'd1873: data <= 8'hF0;
            14'd1874: data <= 8'h00;
            14'd1875: data <= 8'h00;
            14'd1876: data <= 8'h00;
            14'd1877: data <= 8'h00;
            14'd1878: data <= 8'h00;
            14'd1879: data <= 8'h00;
            14'd1880: data <= 8'h00;
            14'd1881: data <= 8'h00;
            14'd1882: data <= 8'h00;
            14'd1883: data <= 8'h00;
            14'd1884: data <= 8'h00;
            14'd1885: data <= 8'h00;
            14'd1886: data <= 8'h0F;
            14'd1887: data <= 8'hFF;
            14'd1888: data <= 8'hFF;
            14'd1889: data <= 8'hFF;
            14'd1890: data <= 8'hFF;
            14'd1891: data <= 8'hFF;
            14'd1892: data <= 8'hFF;
            14'd1893: data <= 8'hFF;
            14'd1894: data <= 8'hFF;
            14'd1895: data <= 8'hFF;
            14'd1896: data <= 8'hFF;
            14'd1897: data <= 8'hFF;
            14'd1898: data <= 8'hFF;
            14'd1899: data <= 8'hFF;
            14'd1900: data <= 8'hFF;
            14'd1901: data <= 8'hFF;
            14'd1902: data <= 8'hFF;
            14'd1903: data <= 8'hFF;
            14'd1904: data <= 8'hFF;
            14'd1905: data <= 8'hFF;
            14'd1906: data <= 8'hFF;
            14'd1907: data <= 8'hFF;
            14'd1908: data <= 8'hFF;
            14'd1909: data <= 8'hFF;
            14'd1910: data <= 8'hFF;
            14'd1911: data <= 8'hFF;
            14'd1912: data <= 8'hFF;
            14'd1913: data <= 8'hF0;
            14'd1914: data <= 8'h00;
            14'd1915: data <= 8'h00;
            14'd1916: data <= 8'h00;
            14'd1917: data <= 8'h00;
            14'd1918: data <= 8'h00;
            14'd1919: data <= 8'h00;
            14'd1920: data <= 8'h00;
            14'd1921: data <= 8'h00;
            14'd1922: data <= 8'h00;
            14'd1923: data <= 8'h00;
            14'd1924: data <= 8'h00;
            14'd1925: data <= 8'h00;
            14'd1926: data <= 8'h0F;
            14'd1927: data <= 8'hFF;
            14'd1928: data <= 8'hFF;
            14'd1929: data <= 8'hFF;
            14'd1930: data <= 8'hFF;
            14'd1931: data <= 8'hFF;
            14'd1932: data <= 8'hFF;
            14'd1933: data <= 8'hFF;
            14'd1934: data <= 8'hFF;
            14'd1935: data <= 8'hFF;
            14'd1936: data <= 8'hFF;
            14'd1937: data <= 8'hFF;
            14'd1938: data <= 8'hFF;
            14'd1939: data <= 8'hFF;
            14'd1940: data <= 8'hFF;
            14'd1941: data <= 8'hFF;
            14'd1942: data <= 8'hFF;
            14'd1943: data <= 8'hFF;
            14'd1944: data <= 8'hFF;
            14'd1945: data <= 8'hFF;
            14'd1946: data <= 8'hFF;
            14'd1947: data <= 8'hFF;
            14'd1948: data <= 8'hFF;
            14'd1949: data <= 8'hFF;
            14'd1950: data <= 8'hFF;
            14'd1951: data <= 8'hFF;
            14'd1952: data <= 8'hFF;
            14'd1953: data <= 8'hF0;
            14'd1954: data <= 8'h00;
            14'd1955: data <= 8'h00;
            14'd1956: data <= 8'h00;
            14'd1957: data <= 8'h00;
            14'd1958: data <= 8'h00;
            14'd1959: data <= 8'h00;
            14'd1960: data <= 8'h00;
            14'd1961: data <= 8'h00;
            14'd1962: data <= 8'h00;
            14'd1963: data <= 8'h00;
            14'd1964: data <= 8'h00;
            14'd1965: data <= 8'h00;
            14'd1966: data <= 8'h0F;
            14'd1967: data <= 8'hFF;
            14'd1968: data <= 8'hFF;
            14'd1969: data <= 8'hFF;
            14'd1970: data <= 8'hFF;
            14'd1971: data <= 8'hFF;
            14'd1972: data <= 8'hFF;
            14'd1973: data <= 8'hFF;
            14'd1974: data <= 8'hFF;
            14'd1975: data <= 8'hFF;
            14'd1976: data <= 8'hFF;
            14'd1977: data <= 8'hFF;
            14'd1978: data <= 8'hFF;
            14'd1979: data <= 8'hFF;
            14'd1980: data <= 8'hFF;
            14'd1981: data <= 8'hFF;
            14'd1982: data <= 8'hFF;
            14'd1983: data <= 8'hFF;
            14'd1984: data <= 8'hFF;
            14'd1985: data <= 8'hFF;
            14'd1986: data <= 8'hFF;
            14'd1987: data <= 8'hFF;
            14'd1988: data <= 8'hFF;
            14'd1989: data <= 8'hFF;
            14'd1990: data <= 8'hFF;
            14'd1991: data <= 8'hFF;
            14'd1992: data <= 8'hFF;
            14'd1993: data <= 8'hF0;
            14'd1994: data <= 8'h00;
            14'd1995: data <= 8'h00;
            14'd1996: data <= 8'h00;
            14'd1997: data <= 8'h00;
            14'd1998: data <= 8'h00;
            14'd1999: data <= 8'h00;
            14'd2000: data <= 8'h00;
            14'd2001: data <= 8'h00;
            14'd2002: data <= 8'h00;
            14'd2003: data <= 8'h00;
            14'd2004: data <= 8'h00;
            14'd2005: data <= 8'h00;
            14'd2006: data <= 8'h0F;
            14'd2007: data <= 8'hFF;
            14'd2008: data <= 8'hFF;
            14'd2009: data <= 8'hFF;
            14'd2010: data <= 8'hFF;
            14'd2011: data <= 8'hFF;
            14'd2012: data <= 8'hFF;
            14'd2013: data <= 8'hFF;
            14'd2014: data <= 8'hFF;
            14'd2015: data <= 8'hFF;
            14'd2016: data <= 8'hFF;
            14'd2017: data <= 8'hFF;
            14'd2018: data <= 8'hFF;
            14'd2019: data <= 8'hFF;
            14'd2020: data <= 8'hFF;
            14'd2021: data <= 8'hFF;
            14'd2022: data <= 8'hFF;
            14'd2023: data <= 8'hFF;
            14'd2024: data <= 8'hFF;
            14'd2025: data <= 8'hFF;
            14'd2026: data <= 8'hFF;
            14'd2027: data <= 8'hFF;
            14'd2028: data <= 8'hFF;
            14'd2029: data <= 8'hFF;
            14'd2030: data <= 8'hFF;
            14'd2031: data <= 8'hFF;
            14'd2032: data <= 8'hFF;
            14'd2033: data <= 8'hF0;
            14'd2034: data <= 8'h00;
            14'd2035: data <= 8'h00;
            14'd2036: data <= 8'h00;
            14'd2037: data <= 8'h00;
            14'd2038: data <= 8'h00;
            14'd2039: data <= 8'h00;
            14'd2040: data <= 8'h00;
            14'd2041: data <= 8'h00;
            14'd2042: data <= 8'h00;
            14'd2043: data <= 8'h00;
            14'd2044: data <= 8'h00;
            14'd2045: data <= 8'h00;
            14'd2046: data <= 8'h0F;
            14'd2047: data <= 8'hFF;
            14'd2048: data <= 8'hFF;
            14'd2049: data <= 8'hFF;
            14'd2050: data <= 8'hFF;
            14'd2051: data <= 8'hFF;
            14'd2052: data <= 8'hFF;
            14'd2053: data <= 8'hFF;
            14'd2054: data <= 8'hFF;
            14'd2055: data <= 8'hFF;
            14'd2056: data <= 8'hFF;
            14'd2057: data <= 8'hFF;
            14'd2058: data <= 8'hFF;
            14'd2059: data <= 8'hFF;
            14'd2060: data <= 8'hFF;
            14'd2061: data <= 8'hFF;
            14'd2062: data <= 8'hFF;
            14'd2063: data <= 8'hFF;
            14'd2064: data <= 8'hFF;
            14'd2065: data <= 8'hFF;
            14'd2066: data <= 8'hFF;
            14'd2067: data <= 8'hFF;
            14'd2068: data <= 8'hFF;
            14'd2069: data <= 8'hFF;
            14'd2070: data <= 8'hFF;
            14'd2071: data <= 8'hFF;
            14'd2072: data <= 8'hFF;
            14'd2073: data <= 8'hF0;
            14'd2074: data <= 8'h00;
            14'd2075: data <= 8'h00;
            14'd2076: data <= 8'h00;
            14'd2077: data <= 8'h00;
            14'd2078: data <= 8'h00;
            14'd2079: data <= 8'h00;
            14'd2080: data <= 8'h00;
            14'd2081: data <= 8'h00;
            14'd2082: data <= 8'h00;
            14'd2083: data <= 8'h00;
            14'd2084: data <= 8'h00;
            14'd2085: data <= 8'h00;
            14'd2086: data <= 8'h0F;
            14'd2087: data <= 8'hFF;
            14'd2088: data <= 8'hFF;
            14'd2089: data <= 8'hFF;
            14'd2090: data <= 8'hFF;
            14'd2091: data <= 8'hFF;
            14'd2092: data <= 8'hFF;
            14'd2093: data <= 8'hFF;
            14'd2094: data <= 8'hFF;
            14'd2095: data <= 8'hFF;
            14'd2096: data <= 8'hFF;
            14'd2097: data <= 8'hFF;
            14'd2098: data <= 8'hFF;
            14'd2099: data <= 8'hFF;
            14'd2100: data <= 8'hFF;
            14'd2101: data <= 8'hFF;
            14'd2102: data <= 8'hFF;
            14'd2103: data <= 8'hFF;
            14'd2104: data <= 8'hFF;
            14'd2105: data <= 8'hFF;
            14'd2106: data <= 8'hFF;
            14'd2107: data <= 8'hFF;
            14'd2108: data <= 8'hFF;
            14'd2109: data <= 8'hFF;
            14'd2110: data <= 8'hFF;
            14'd2111: data <= 8'hFF;
            14'd2112: data <= 8'hFF;
            14'd2113: data <= 8'hF0;
            14'd2114: data <= 8'h00;
            14'd2115: data <= 8'h00;
            14'd2116: data <= 8'h00;
            14'd2117: data <= 8'h00;
            14'd2118: data <= 8'h00;
            14'd2119: data <= 8'h00;
            14'd2120: data <= 8'h00;
            14'd2121: data <= 8'h00;
            14'd2122: data <= 8'h00;
            14'd2123: data <= 8'h00;
            14'd2124: data <= 8'h00;
            14'd2125: data <= 8'h00;
            14'd2126: data <= 8'h0F;
            14'd2127: data <= 8'hFF;
            14'd2128: data <= 8'hFF;
            14'd2129: data <= 8'hFF;
            14'd2130: data <= 8'hFF;
            14'd2131: data <= 8'hFF;
            14'd2132: data <= 8'hFF;
            14'd2133: data <= 8'hFF;
            14'd2134: data <= 8'hFF;
            14'd2135: data <= 8'hFF;
            14'd2136: data <= 8'hFF;
            14'd2137: data <= 8'hFF;
            14'd2138: data <= 8'hFF;
            14'd2139: data <= 8'hFF;
            14'd2140: data <= 8'hFF;
            14'd2141: data <= 8'hFF;
            14'd2142: data <= 8'hFF;
            14'd2143: data <= 8'hFF;
            14'd2144: data <= 8'hFF;
            14'd2145: data <= 8'hFF;
            14'd2146: data <= 8'hFF;
            14'd2147: data <= 8'hFF;
            14'd2148: data <= 8'hFF;
            14'd2149: data <= 8'hFF;
            14'd2150: data <= 8'hFF;
            14'd2151: data <= 8'hFF;
            14'd2152: data <= 8'hFF;
            14'd2153: data <= 8'hF0;
            14'd2154: data <= 8'h00;
            14'd2155: data <= 8'h00;
            14'd2156: data <= 8'h00;
            14'd2157: data <= 8'h00;
            14'd2158: data <= 8'h00;
            14'd2159: data <= 8'h00;
            14'd2160: data <= 8'h00;
            14'd2161: data <= 8'h00;
            14'd2162: data <= 8'h00;
            14'd2163: data <= 8'h00;
            14'd2164: data <= 8'h00;
            14'd2165: data <= 8'h00;
            14'd2166: data <= 8'h0F;
            14'd2167: data <= 8'hFF;
            14'd2168: data <= 8'hFF;
            14'd2169: data <= 8'hFF;
            14'd2170: data <= 8'hFF;
            14'd2171: data <= 8'hFF;
            14'd2172: data <= 8'hFF;
            14'd2173: data <= 8'hFF;
            14'd2174: data <= 8'hFF;
            14'd2175: data <= 8'hFF;
            14'd2176: data <= 8'hFF;
            14'd2177: data <= 8'hFF;
            14'd2178: data <= 8'hFF;
            14'd2179: data <= 8'hFF;
            14'd2180: data <= 8'hFF;
            14'd2181: data <= 8'hFF;
            14'd2182: data <= 8'hFF;
            14'd2183: data <= 8'hFF;
            14'd2184: data <= 8'hFF;
            14'd2185: data <= 8'hFF;
            14'd2186: data <= 8'hFF;
            14'd2187: data <= 8'hFF;
            14'd2188: data <= 8'hFF;
            14'd2189: data <= 8'hFF;
            14'd2190: data <= 8'hFF;
            14'd2191: data <= 8'hFF;
            14'd2192: data <= 8'hFF;
            14'd2193: data <= 8'hF0;
            14'd2194: data <= 8'h00;
            14'd2195: data <= 8'h00;
            14'd2196: data <= 8'h00;
            14'd2197: data <= 8'h00;
            14'd2198: data <= 8'h00;
            14'd2199: data <= 8'h00;
            14'd2200: data <= 8'h00;
            14'd2201: data <= 8'h00;
            14'd2202: data <= 8'h00;
            14'd2203: data <= 8'h00;
            14'd2204: data <= 8'h00;
            14'd2205: data <= 8'h00;
            14'd2206: data <= 8'h0F;
            14'd2207: data <= 8'hFF;
            14'd2208: data <= 8'hFF;
            14'd2209: data <= 8'hFF;
            14'd2210: data <= 8'hFF;
            14'd2211: data <= 8'hFF;
            14'd2212: data <= 8'hFF;
            14'd2213: data <= 8'hFF;
            14'd2214: data <= 8'hFF;
            14'd2215: data <= 8'hFF;
            14'd2216: data <= 8'hFF;
            14'd2217: data <= 8'hFD;
            14'd2218: data <= 8'hFF;
            14'd2219: data <= 8'hFF;
            14'd2220: data <= 8'hFF;
            14'd2221: data <= 8'hFF;
            14'd2222: data <= 8'hFF;
            14'd2223: data <= 8'hFF;
            14'd2224: data <= 8'hFF;
            14'd2225: data <= 8'hFF;
            14'd2226: data <= 8'hFF;
            14'd2227: data <= 8'hFF;
            14'd2228: data <= 8'hFF;
            14'd2229: data <= 8'hFF;
            14'd2230: data <= 8'hFF;
            14'd2231: data <= 8'hFF;
            14'd2232: data <= 8'hFF;
            14'd2233: data <= 8'hF0;
            14'd2234: data <= 8'h00;
            14'd2235: data <= 8'h00;
            14'd2236: data <= 8'h00;
            14'd2237: data <= 8'h00;
            14'd2238: data <= 8'h00;
            14'd2239: data <= 8'h00;
            14'd2240: data <= 8'h00;
            14'd2241: data <= 8'h00;
            14'd2242: data <= 8'h00;
            14'd2243: data <= 8'h00;
            14'd2244: data <= 8'h00;
            14'd2245: data <= 8'h00;
            14'd2246: data <= 8'h0F;
            14'd2247: data <= 8'hFF;
            14'd2248: data <= 8'hFF;
            14'd2249: data <= 8'hFF;
            14'd2250: data <= 8'hFF;
            14'd2251: data <= 8'hFF;
            14'd2252: data <= 8'hFF;
            14'd2253: data <= 8'hFF;
            14'd2254: data <= 8'hFF;
            14'd2255: data <= 8'hFF;
            14'd2256: data <= 8'hFF;
            14'd2257: data <= 8'hFF;
            14'd2258: data <= 8'hFF;
            14'd2259: data <= 8'hFF;
            14'd2260: data <= 8'hFF;
            14'd2261: data <= 8'hFF;
            14'd2262: data <= 8'hFF;
            14'd2263: data <= 8'hFF;
            14'd2264: data <= 8'hFF;
            14'd2265: data <= 8'hFF;
            14'd2266: data <= 8'hFF;
            14'd2267: data <= 8'hFF;
            14'd2268: data <= 8'hFF;
            14'd2269: data <= 8'hFF;
            14'd2270: data <= 8'hFF;
            14'd2271: data <= 8'hFF;
            14'd2272: data <= 8'hFF;
            14'd2273: data <= 8'hF0;
            14'd2274: data <= 8'h00;
            14'd2275: data <= 8'h00;
            14'd2276: data <= 8'h00;
            14'd2277: data <= 8'h00;
            14'd2278: data <= 8'h00;
            14'd2279: data <= 8'h00;
            14'd2280: data <= 8'h00;
            14'd2281: data <= 8'h00;
            14'd2282: data <= 8'h00;
            14'd2283: data <= 8'h00;
            14'd2284: data <= 8'h00;
            14'd2285: data <= 8'h00;
            14'd2286: data <= 8'h0F;
            14'd2287: data <= 8'hFF;
            14'd2288: data <= 8'hFF;
            14'd2289: data <= 8'hFF;
            14'd2290: data <= 8'hFF;
            14'd2291: data <= 8'hFF;
            14'd2292: data <= 8'hFF;
            14'd2293: data <= 8'hFF;
            14'd2294: data <= 8'hFF;
            14'd2295: data <= 8'hFF;
            14'd2296: data <= 8'hFF;
            14'd2297: data <= 8'hFF;
            14'd2298: data <= 8'hFF;
            14'd2299: data <= 8'hFF;
            14'd2300: data <= 8'hFF;
            14'd2301: data <= 8'hFF;
            14'd2302: data <= 8'hFF;
            14'd2303: data <= 8'hFF;
            14'd2304: data <= 8'hFF;
            14'd2305: data <= 8'hFF;
            14'd2306: data <= 8'hFF;
            14'd2307: data <= 8'hFF;
            14'd2308: data <= 8'hFF;
            14'd2309: data <= 8'hFF;
            14'd2310: data <= 8'hFF;
            14'd2311: data <= 8'hFF;
            14'd2312: data <= 8'hFF;
            14'd2313: data <= 8'hF0;
            14'd2314: data <= 8'h00;
            14'd2315: data <= 8'h00;
            14'd2316: data <= 8'h00;
            14'd2317: data <= 8'h00;
            14'd2318: data <= 8'h00;
            14'd2319: data <= 8'h00;
            14'd2320: data <= 8'h00;
            14'd2321: data <= 8'h00;
            14'd2322: data <= 8'h00;
            14'd2323: data <= 8'h00;
            14'd2324: data <= 8'h00;
            14'd2325: data <= 8'h00;
            14'd2326: data <= 8'h0F;
            14'd2327: data <= 8'hFF;
            14'd2328: data <= 8'hFF;
            14'd2329: data <= 8'hFF;
            14'd2330: data <= 8'hFF;
            14'd2331: data <= 8'hFF;
            14'd2332: data <= 8'hFF;
            14'd2333: data <= 8'hFF;
            14'd2334: data <= 8'hFF;
            14'd2335: data <= 8'hFF;
            14'd2336: data <= 8'hFF;
            14'd2337: data <= 8'hFF;
            14'd2338: data <= 8'hFF;
            14'd2339: data <= 8'hFF;
            14'd2340: data <= 8'hFF;
            14'd2341: data <= 8'hFF;
            14'd2342: data <= 8'hFF;
            14'd2343: data <= 8'hFF;
            14'd2344: data <= 8'hFF;
            14'd2345: data <= 8'hFF;
            14'd2346: data <= 8'hFF;
            14'd2347: data <= 8'hFF;
            14'd2348: data <= 8'hF7;
            14'd2349: data <= 8'hFF;
            14'd2350: data <= 8'hFF;
            14'd2351: data <= 8'hFF;
            14'd2352: data <= 8'hFF;
            14'd2353: data <= 8'hF0;
            14'd2354: data <= 8'h00;
            14'd2355: data <= 8'h00;
            14'd2356: data <= 8'h00;
            14'd2357: data <= 8'h00;
            14'd2358: data <= 8'h00;
            14'd2359: data <= 8'h00;
            14'd2360: data <= 8'h00;
            14'd2361: data <= 8'h00;
            14'd2362: data <= 8'h00;
            14'd2363: data <= 8'h00;
            14'd2364: data <= 8'h00;
            14'd2365: data <= 8'h00;
            14'd2366: data <= 8'h0F;
            14'd2367: data <= 8'hFF;
            14'd2368: data <= 8'hFF;
            14'd2369: data <= 8'hFF;
            14'd2370: data <= 8'hFF;
            14'd2371: data <= 8'hFF;
            14'd2372: data <= 8'hFF;
            14'd2373: data <= 8'hFF;
            14'd2374: data <= 8'hFF;
            14'd2375: data <= 8'hFF;
            14'd2376: data <= 8'hFF;
            14'd2377: data <= 8'hFF;
            14'd2378: data <= 8'hFF;
            14'd2379: data <= 8'hFF;
            14'd2380: data <= 8'hFF;
            14'd2381: data <= 8'hFF;
            14'd2382: data <= 8'hFF;
            14'd2383: data <= 8'hFF;
            14'd2384: data <= 8'hFF;
            14'd2385: data <= 8'hFF;
            14'd2386: data <= 8'hFF;
            14'd2387: data <= 8'hFF;
            14'd2388: data <= 8'hFF;
            14'd2389: data <= 8'hFF;
            14'd2390: data <= 8'hFF;
            14'd2391: data <= 8'hFF;
            14'd2392: data <= 8'hFF;
            14'd2393: data <= 8'hF0;
            14'd2394: data <= 8'h00;
            14'd2395: data <= 8'h00;
            14'd2396: data <= 8'h00;
            14'd2397: data <= 8'h00;
            14'd2398: data <= 8'h00;
            14'd2399: data <= 8'h00;
            14'd2400: data <= 8'h00;
            14'd2401: data <= 8'h00;
            14'd2402: data <= 8'h00;
            14'd2403: data <= 8'h00;
            14'd2404: data <= 8'h00;
            14'd2405: data <= 8'h00;
            14'd2406: data <= 8'h0F;
            14'd2407: data <= 8'hFF;
            14'd2408: data <= 8'hFF;
            14'd2409: data <= 8'hFF;
            14'd2410: data <= 8'hFF;
            14'd2411: data <= 8'hFF;
            14'd2412: data <= 8'hFF;
            14'd2413: data <= 8'hFF;
            14'd2414: data <= 8'hFF;
            14'd2415: data <= 8'hFF;
            14'd2416: data <= 8'hFF;
            14'd2417: data <= 8'hFF;
            14'd2418: data <= 8'hFF;
            14'd2419: data <= 8'hFF;
            14'd2420: data <= 8'hFF;
            14'd2421: data <= 8'hFF;
            14'd2422: data <= 8'hFF;
            14'd2423: data <= 8'hFF;
            14'd2424: data <= 8'hFF;
            14'd2425: data <= 8'hFF;
            14'd2426: data <= 8'hFF;
            14'd2427: data <= 8'hFF;
            14'd2428: data <= 8'hFF;
            14'd2429: data <= 8'hFF;
            14'd2430: data <= 8'hFF;
            14'd2431: data <= 8'hFF;
            14'd2432: data <= 8'hFF;
            14'd2433: data <= 8'hF0;
            14'd2434: data <= 8'h00;
            14'd2435: data <= 8'h00;
            14'd2436: data <= 8'h00;
            14'd2437: data <= 8'h00;
            14'd2438: data <= 8'h00;
            14'd2439: data <= 8'h00;
            14'd2440: data <= 8'h00;
            14'd2441: data <= 8'h00;
            14'd2442: data <= 8'h00;
            14'd2443: data <= 8'h00;
            14'd2444: data <= 8'h00;
            14'd2445: data <= 8'h00;
            14'd2446: data <= 8'h0F;
            14'd2447: data <= 8'hFF;
            14'd2448: data <= 8'hFF;
            14'd2449: data <= 8'hFF;
            14'd2450: data <= 8'hFF;
            14'd2451: data <= 8'hFF;
            14'd2452: data <= 8'hFF;
            14'd2453: data <= 8'hFF;
            14'd2454: data <= 8'hFF;
            14'd2455: data <= 8'hFF;
            14'd2456: data <= 8'hFF;
            14'd2457: data <= 8'hFF;
            14'd2458: data <= 8'hFF;
            14'd2459: data <= 8'hFF;
            14'd2460: data <= 8'hFF;
            14'd2461: data <= 8'hFF;
            14'd2462: data <= 8'hFF;
            14'd2463: data <= 8'hFF;
            14'd2464: data <= 8'hFF;
            14'd2465: data <= 8'hFF;
            14'd2466: data <= 8'hFF;
            14'd2467: data <= 8'hFF;
            14'd2468: data <= 8'hFF;
            14'd2469: data <= 8'hFF;
            14'd2470: data <= 8'hFF;
            14'd2471: data <= 8'hFF;
            14'd2472: data <= 8'hFF;
            14'd2473: data <= 8'hF0;
            14'd2474: data <= 8'h00;
            14'd2475: data <= 8'h00;
            14'd2476: data <= 8'h00;
            14'd2477: data <= 8'h00;
            14'd2478: data <= 8'h00;
            14'd2479: data <= 8'h00;
            14'd2480: data <= 8'h00;
            14'd2481: data <= 8'h00;
            14'd2482: data <= 8'h00;
            14'd2483: data <= 8'h00;
            14'd2484: data <= 8'h00;
            14'd2485: data <= 8'h00;
            14'd2486: data <= 8'h0F;
            14'd2487: data <= 8'hFF;
            14'd2488: data <= 8'hFF;
            14'd2489: data <= 8'hFF;
            14'd2490: data <= 8'hFF;
            14'd2491: data <= 8'hFF;
            14'd2492: data <= 8'hFF;
            14'd2493: data <= 8'hFF;
            14'd2494: data <= 8'hFF;
            14'd2495: data <= 8'hFF;
            14'd2496: data <= 8'hE7;
            14'd2497: data <= 8'hFF;
            14'd2498: data <= 8'hFF;
            14'd2499: data <= 8'hFF;
            14'd2500: data <= 8'hFF;
            14'd2501: data <= 8'hFF;
            14'd2502: data <= 8'hFF;
            14'd2503: data <= 8'h0F;
            14'd2504: data <= 8'hFF;
            14'd2505: data <= 8'hFF;
            14'd2506: data <= 8'hFF;
            14'd2507: data <= 8'hFF;
            14'd2508: data <= 8'hFF;
            14'd2509: data <= 8'hFF;
            14'd2510: data <= 8'hFF;
            14'd2511: data <= 8'hFF;
            14'd2512: data <= 8'hFF;
            14'd2513: data <= 8'hF0;
            14'd2514: data <= 8'h00;
            14'd2515: data <= 8'h00;
            14'd2516: data <= 8'h00;
            14'd2517: data <= 8'h00;
            14'd2518: data <= 8'h00;
            14'd2519: data <= 8'h00;
            14'd2520: data <= 8'h00;
            14'd2521: data <= 8'h00;
            14'd2522: data <= 8'h00;
            14'd2523: data <= 8'h00;
            14'd2524: data <= 8'h00;
            14'd2525: data <= 8'h00;
            14'd2526: data <= 8'h0F;
            14'd2527: data <= 8'hFF;
            14'd2528: data <= 8'hFF;
            14'd2529: data <= 8'hFF;
            14'd2530: data <= 8'hFF;
            14'd2531: data <= 8'hFF;
            14'd2532: data <= 8'hFF;
            14'd2533: data <= 8'hFF;
            14'd2534: data <= 8'hFF;
            14'd2535: data <= 8'hFF;
            14'd2536: data <= 8'h80;
            14'd2537: data <= 8'hFF;
            14'd2538: data <= 8'hFF;
            14'd2539: data <= 8'hFF;
            14'd2540: data <= 8'hFF;
            14'd2541: data <= 8'hFF;
            14'd2542: data <= 8'hFC;
            14'd2543: data <= 8'h07;
            14'd2544: data <= 8'hFD;
            14'd2545: data <= 8'hFF;
            14'd2546: data <= 8'hFF;
            14'd2547: data <= 8'hFF;
            14'd2548: data <= 8'hFF;
            14'd2549: data <= 8'hFF;
            14'd2550: data <= 8'hFF;
            14'd2551: data <= 8'hFF;
            14'd2552: data <= 8'hFF;
            14'd2553: data <= 8'hF0;
            14'd2554: data <= 8'h00;
            14'd2555: data <= 8'h00;
            14'd2556: data <= 8'h00;
            14'd2557: data <= 8'h00;
            14'd2558: data <= 8'h00;
            14'd2559: data <= 8'h00;
            14'd2560: data <= 8'h00;
            14'd2561: data <= 8'h00;
            14'd2562: data <= 8'h00;
            14'd2563: data <= 8'h00;
            14'd2564: data <= 8'h00;
            14'd2565: data <= 8'h00;
            14'd2566: data <= 8'h0F;
            14'd2567: data <= 8'hFF;
            14'd2568: data <= 8'hFF;
            14'd2569: data <= 8'hFF;
            14'd2570: data <= 8'hFF;
            14'd2571: data <= 8'hFF;
            14'd2572: data <= 8'hFF;
            14'd2573: data <= 8'hFF;
            14'd2574: data <= 8'hFF;
            14'd2575: data <= 8'hFF;
            14'd2576: data <= 8'h80;
            14'd2577: data <= 8'h1F;
            14'd2578: data <= 8'hFF;
            14'd2579: data <= 8'hFF;
            14'd2580: data <= 8'hFF;
            14'd2581: data <= 8'hFF;
            14'd2582: data <= 8'hF0;
            14'd2583: data <= 8'h03;
            14'd2584: data <= 8'hFF;
            14'd2585: data <= 8'hFF;
            14'd2586: data <= 8'hFF;
            14'd2587: data <= 8'hFF;
            14'd2588: data <= 8'hFF;
            14'd2589: data <= 8'hFF;
            14'd2590: data <= 8'hFF;
            14'd2591: data <= 8'hFF;
            14'd2592: data <= 8'hFF;
            14'd2593: data <= 8'hF0;
            14'd2594: data <= 8'h00;
            14'd2595: data <= 8'h00;
            14'd2596: data <= 8'h00;
            14'd2597: data <= 8'h00;
            14'd2598: data <= 8'h00;
            14'd2599: data <= 8'h00;
            14'd2600: data <= 8'h00;
            14'd2601: data <= 8'h00;
            14'd2602: data <= 8'h00;
            14'd2603: data <= 8'h00;
            14'd2604: data <= 8'h00;
            14'd2605: data <= 8'h00;
            14'd2606: data <= 8'h0F;
            14'd2607: data <= 8'hFF;
            14'd2608: data <= 8'hFF;
            14'd2609: data <= 8'hFF;
            14'd2610: data <= 8'hFF;
            14'd2611: data <= 8'hFF;
            14'd2612: data <= 8'hFF;
            14'd2613: data <= 8'hFF;
            14'd2614: data <= 8'hFF;
            14'd2615: data <= 8'hFF;
            14'd2616: data <= 8'h00;
            14'd2617: data <= 8'h01;
            14'd2618: data <= 8'hFF;
            14'd2619: data <= 8'hFF;
            14'd2620: data <= 8'hFF;
            14'd2621: data <= 8'hFF;
            14'd2622: data <= 8'hC0;
            14'd2623: data <= 8'h07;
            14'd2624: data <= 8'hFF;
            14'd2625: data <= 8'hFF;
            14'd2626: data <= 8'hFF;
            14'd2627: data <= 8'hFF;
            14'd2628: data <= 8'hFF;
            14'd2629: data <= 8'hFF;
            14'd2630: data <= 8'hFF;
            14'd2631: data <= 8'hFF;
            14'd2632: data <= 8'hFF;
            14'd2633: data <= 8'hF0;
            14'd2634: data <= 8'h00;
            14'd2635: data <= 8'h00;
            14'd2636: data <= 8'h00;
            14'd2637: data <= 8'h00;
            14'd2638: data <= 8'h00;
            14'd2639: data <= 8'h00;
            14'd2640: data <= 8'h00;
            14'd2641: data <= 8'h00;
            14'd2642: data <= 8'h00;
            14'd2643: data <= 8'h00;
            14'd2644: data <= 8'h00;
            14'd2645: data <= 8'h00;
            14'd2646: data <= 8'h0F;
            14'd2647: data <= 8'hFF;
            14'd2648: data <= 8'hFF;
            14'd2649: data <= 8'hFF;
            14'd2650: data <= 8'hFF;
            14'd2651: data <= 8'hFF;
            14'd2652: data <= 8'hFF;
            14'd2653: data <= 8'hFF;
            14'd2654: data <= 8'hFF;
            14'd2655: data <= 8'hFF;
            14'd2656: data <= 8'h80;
            14'd2657: data <= 8'h00;
            14'd2658: data <= 8'h3F;
            14'd2659: data <= 8'hFF;
            14'd2660: data <= 8'hFF;
            14'd2661: data <= 8'hFF;
            14'd2662: data <= 8'h80;
            14'd2663: data <= 8'h07;
            14'd2664: data <= 8'hFF;
            14'd2665: data <= 8'hFF;
            14'd2666: data <= 8'hFF;
            14'd2667: data <= 8'hFF;
            14'd2668: data <= 8'hFF;
            14'd2669: data <= 8'hFF;
            14'd2670: data <= 8'hFF;
            14'd2671: data <= 8'hFF;
            14'd2672: data <= 8'hFF;
            14'd2673: data <= 8'hF0;
            14'd2674: data <= 8'h00;
            14'd2675: data <= 8'h00;
            14'd2676: data <= 8'h00;
            14'd2677: data <= 8'h00;
            14'd2678: data <= 8'h00;
            14'd2679: data <= 8'h00;
            14'd2680: data <= 8'h00;
            14'd2681: data <= 8'h00;
            14'd2682: data <= 8'h00;
            14'd2683: data <= 8'h00;
            14'd2684: data <= 8'h00;
            14'd2685: data <= 8'h00;
            14'd2686: data <= 8'h0F;
            14'd2687: data <= 8'hFF;
            14'd2688: data <= 8'hFF;
            14'd2689: data <= 8'hFF;
            14'd2690: data <= 8'hFF;
            14'd2691: data <= 8'hFF;
            14'd2692: data <= 8'hFF;
            14'd2693: data <= 8'hFF;
            14'd2694: data <= 8'hFF;
            14'd2695: data <= 8'hFD;
            14'd2696: data <= 8'h80;
            14'd2697: data <= 8'h00;
            14'd2698: data <= 8'h07;
            14'd2699: data <= 8'hFF;
            14'd2700: data <= 8'hFF;
            14'd2701: data <= 8'hFE;
            14'd2702: data <= 8'h00;
            14'd2703: data <= 8'h0F;
            14'd2704: data <= 8'hFF;
            14'd2705: data <= 8'hFF;
            14'd2706: data <= 8'hFF;
            14'd2707: data <= 8'hFF;
            14'd2708: data <= 8'hFF;
            14'd2709: data <= 8'hFF;
            14'd2710: data <= 8'hFF;
            14'd2711: data <= 8'hFF;
            14'd2712: data <= 8'hFF;
            14'd2713: data <= 8'hF0;
            14'd2714: data <= 8'h00;
            14'd2715: data <= 8'h00;
            14'd2716: data <= 8'h00;
            14'd2717: data <= 8'h00;
            14'd2718: data <= 8'h00;
            14'd2719: data <= 8'h00;
            14'd2720: data <= 8'h00;
            14'd2721: data <= 8'h00;
            14'd2722: data <= 8'h00;
            14'd2723: data <= 8'h00;
            14'd2724: data <= 8'h00;
            14'd2725: data <= 8'h00;
            14'd2726: data <= 8'h0F;
            14'd2727: data <= 8'hFF;
            14'd2728: data <= 8'hFF;
            14'd2729: data <= 8'hFF;
            14'd2730: data <= 8'hFF;
            14'd2731: data <= 8'hFF;
            14'd2732: data <= 8'hFF;
            14'd2733: data <= 8'hFF;
            14'd2734: data <= 8'hFF;
            14'd2735: data <= 8'hFF;
            14'd2736: data <= 8'hF0;
            14'd2737: data <= 8'h00;
            14'd2738: data <= 8'h07;
            14'd2739: data <= 8'hFF;
            14'd2740: data <= 8'hFF;
            14'd2741: data <= 8'hF8;
            14'd2742: data <= 8'h00;
            14'd2743: data <= 8'h7F;
            14'd2744: data <= 8'hFF;
            14'd2745: data <= 8'hFF;
            14'd2746: data <= 8'hFF;
            14'd2747: data <= 8'hFF;
            14'd2748: data <= 8'hFF;
            14'd2749: data <= 8'hFF;
            14'd2750: data <= 8'hFF;
            14'd2751: data <= 8'hFF;
            14'd2752: data <= 8'hFF;
            14'd2753: data <= 8'hF0;
            14'd2754: data <= 8'h00;
            14'd2755: data <= 8'h00;
            14'd2756: data <= 8'h00;
            14'd2757: data <= 8'h00;
            14'd2758: data <= 8'h00;
            14'd2759: data <= 8'h00;
            14'd2760: data <= 8'h00;
            14'd2761: data <= 8'h00;
            14'd2762: data <= 8'h00;
            14'd2763: data <= 8'h00;
            14'd2764: data <= 8'h00;
            14'd2765: data <= 8'h00;
            14'd2766: data <= 8'h0F;
            14'd2767: data <= 8'hFF;
            14'd2768: data <= 8'hFF;
            14'd2769: data <= 8'hFF;
            14'd2770: data <= 8'hFF;
            14'd2771: data <= 8'hFF;
            14'd2772: data <= 8'hFF;
            14'd2773: data <= 8'hFF;
            14'd2774: data <= 8'hFF;
            14'd2775: data <= 8'hFF;
            14'd2776: data <= 8'hFE;
            14'd2777: data <= 8'h00;
            14'd2778: data <= 8'h03;
            14'd2779: data <= 8'hFF;
            14'd2780: data <= 8'h7F;
            14'd2781: data <= 8'hF0;
            14'd2782: data <= 8'h01;
            14'd2783: data <= 8'hFF;
            14'd2784: data <= 8'hFF;
            14'd2785: data <= 8'hFF;
            14'd2786: data <= 8'hFF;
            14'd2787: data <= 8'hFF;
            14'd2788: data <= 8'hFF;
            14'd2789: data <= 8'hFF;
            14'd2790: data <= 8'hFF;
            14'd2791: data <= 8'hFF;
            14'd2792: data <= 8'hFF;
            14'd2793: data <= 8'hF0;
            14'd2794: data <= 8'h00;
            14'd2795: data <= 8'h00;
            14'd2796: data <= 8'h00;
            14'd2797: data <= 8'h00;
            14'd2798: data <= 8'h00;
            14'd2799: data <= 8'h00;
            14'd2800: data <= 8'h00;
            14'd2801: data <= 8'h00;
            14'd2802: data <= 8'h00;
            14'd2803: data <= 8'h00;
            14'd2804: data <= 8'h00;
            14'd2805: data <= 8'h00;
            14'd2806: data <= 8'h0F;
            14'd2807: data <= 8'hFF;
            14'd2808: data <= 8'hFF;
            14'd2809: data <= 8'hFF;
            14'd2810: data <= 8'hFF;
            14'd2811: data <= 8'hFF;
            14'd2812: data <= 8'hFF;
            14'd2813: data <= 8'hFF;
            14'd2814: data <= 8'hFF;
            14'd2815: data <= 8'hFF;
            14'd2816: data <= 8'hFF;
            14'd2817: data <= 8'h00;
            14'd2818: data <= 8'h03;
            14'd2819: data <= 8'hFF;
            14'd2820: data <= 8'hFF;
            14'd2821: data <= 8'hE0;
            14'd2822: data <= 8'h07;
            14'd2823: data <= 8'hFF;
            14'd2824: data <= 8'hFF;
            14'd2825: data <= 8'hFF;
            14'd2826: data <= 8'hFF;
            14'd2827: data <= 8'hFF;
            14'd2828: data <= 8'hFF;
            14'd2829: data <= 8'hFF;
            14'd2830: data <= 8'hFF;
            14'd2831: data <= 8'hFF;
            14'd2832: data <= 8'hFF;
            14'd2833: data <= 8'hF0;
            14'd2834: data <= 8'h00;
            14'd2835: data <= 8'h00;
            14'd2836: data <= 8'h00;
            14'd2837: data <= 8'h00;
            14'd2838: data <= 8'h00;
            14'd2839: data <= 8'h00;
            14'd2840: data <= 8'h00;
            14'd2841: data <= 8'h00;
            14'd2842: data <= 8'h00;
            14'd2843: data <= 8'h00;
            14'd2844: data <= 8'h00;
            14'd2845: data <= 8'h00;
            14'd2846: data <= 8'h0F;
            14'd2847: data <= 8'hFF;
            14'd2848: data <= 8'hFF;
            14'd2849: data <= 8'hFF;
            14'd2850: data <= 8'hFF;
            14'd2851: data <= 8'hFF;
            14'd2852: data <= 8'hFF;
            14'd2853: data <= 8'hFF;
            14'd2854: data <= 8'hFF;
            14'd2855: data <= 8'hFF;
            14'd2856: data <= 8'hFF;
            14'd2857: data <= 8'hE0;
            14'd2858: data <= 8'h07;
            14'd2859: data <= 8'hFF;
            14'd2860: data <= 8'hFF;
            14'd2861: data <= 8'hC0;
            14'd2862: data <= 8'h0F;
            14'd2863: data <= 8'hFF;
            14'd2864: data <= 8'hFF;
            14'd2865: data <= 8'hFF;
            14'd2866: data <= 8'hFF;
            14'd2867: data <= 8'hFF;
            14'd2868: data <= 8'hFF;
            14'd2869: data <= 8'hFF;
            14'd2870: data <= 8'hFF;
            14'd2871: data <= 8'hFF;
            14'd2872: data <= 8'hFF;
            14'd2873: data <= 8'hF0;
            14'd2874: data <= 8'h00;
            14'd2875: data <= 8'h00;
            14'd2876: data <= 8'h00;
            14'd2877: data <= 8'h00;
            14'd2878: data <= 8'h00;
            14'd2879: data <= 8'h00;
            14'd2880: data <= 8'h00;
            14'd2881: data <= 8'h00;
            14'd2882: data <= 8'h00;
            14'd2883: data <= 8'h00;
            14'd2884: data <= 8'h00;
            14'd2885: data <= 8'h00;
            14'd2886: data <= 8'h0F;
            14'd2887: data <= 8'hFF;
            14'd2888: data <= 8'hFF;
            14'd2889: data <= 8'hFF;
            14'd2890: data <= 8'hFF;
            14'd2891: data <= 8'hFF;
            14'd2892: data <= 8'hFF;
            14'd2893: data <= 8'hFF;
            14'd2894: data <= 8'hFF;
            14'd2895: data <= 8'hFF;
            14'd2896: data <= 8'hFF;
            14'd2897: data <= 8'hFE;
            14'd2898: data <= 8'h0F;
            14'd2899: data <= 8'hFF;
            14'd2900: data <= 8'hFF;
            14'd2901: data <= 8'hC0;
            14'd2902: data <= 8'h3F;
            14'd2903: data <= 8'hFF;
            14'd2904: data <= 8'hFF;
            14'd2905: data <= 8'hFF;
            14'd2906: data <= 8'hFF;
            14'd2907: data <= 8'hFF;
            14'd2908: data <= 8'hFF;
            14'd2909: data <= 8'hFF;
            14'd2910: data <= 8'hFF;
            14'd2911: data <= 8'hFF;
            14'd2912: data <= 8'hFF;
            14'd2913: data <= 8'hF0;
            14'd2914: data <= 8'h00;
            14'd2915: data <= 8'h00;
            14'd2916: data <= 8'h00;
            14'd2917: data <= 8'h00;
            14'd2918: data <= 8'h00;
            14'd2919: data <= 8'h00;
            14'd2920: data <= 8'h00;
            14'd2921: data <= 8'h00;
            14'd2922: data <= 8'h00;
            14'd2923: data <= 8'h00;
            14'd2924: data <= 8'h00;
            14'd2925: data <= 8'h00;
            14'd2926: data <= 8'h0F;
            14'd2927: data <= 8'hFF;
            14'd2928: data <= 8'hFF;
            14'd2929: data <= 8'hFF;
            14'd2930: data <= 8'hFF;
            14'd2931: data <= 8'hFF;
            14'd2932: data <= 8'hFF;
            14'd2933: data <= 8'hFF;
            14'd2934: data <= 8'hFF;
            14'd2935: data <= 8'hFF;
            14'd2936: data <= 8'hFF;
            14'd2937: data <= 8'hFF;
            14'd2938: data <= 8'hFF;
            14'd2939: data <= 8'hFF;
            14'd2940: data <= 8'hFF;
            14'd2941: data <= 8'hC0;
            14'd2942: data <= 8'hFF;
            14'd2943: data <= 8'hFF;
            14'd2944: data <= 8'hFF;
            14'd2945: data <= 8'hFF;
            14'd2946: data <= 8'hFF;
            14'd2947: data <= 8'hFF;
            14'd2948: data <= 8'hFF;
            14'd2949: data <= 8'hFF;
            14'd2950: data <= 8'hFF;
            14'd2951: data <= 8'hFF;
            14'd2952: data <= 8'hFF;
            14'd2953: data <= 8'hF0;
            14'd2954: data <= 8'h00;
            14'd2955: data <= 8'h00;
            14'd2956: data <= 8'h00;
            14'd2957: data <= 8'h00;
            14'd2958: data <= 8'h00;
            14'd2959: data <= 8'h00;
            14'd2960: data <= 8'h00;
            14'd2961: data <= 8'h00;
            14'd2962: data <= 8'h00;
            14'd2963: data <= 8'h00;
            14'd2964: data <= 8'h00;
            14'd2965: data <= 8'h00;
            14'd2966: data <= 8'h0F;
            14'd2967: data <= 8'hFF;
            14'd2968: data <= 8'hFF;
            14'd2969: data <= 8'hFF;
            14'd2970: data <= 8'hFF;
            14'd2971: data <= 8'hFF;
            14'd2972: data <= 8'hFF;
            14'd2973: data <= 8'hFF;
            14'd2974: data <= 8'hFF;
            14'd2975: data <= 8'hFF;
            14'd2976: data <= 8'hFF;
            14'd2977: data <= 8'hFF;
            14'd2978: data <= 8'hFF;
            14'd2979: data <= 8'hFF;
            14'd2980: data <= 8'hFF;
            14'd2981: data <= 8'hE3;
            14'd2982: data <= 8'hFF;
            14'd2983: data <= 8'hFF;
            14'd2984: data <= 8'hFF;
            14'd2985: data <= 8'hFF;
            14'd2986: data <= 8'hFF;
            14'd2987: data <= 8'hFF;
            14'd2988: data <= 8'hFF;
            14'd2989: data <= 8'hFF;
            14'd2990: data <= 8'hFF;
            14'd2991: data <= 8'hFF;
            14'd2992: data <= 8'hFF;
            14'd2993: data <= 8'hF0;
            14'd2994: data <= 8'h00;
            14'd2995: data <= 8'h00;
            14'd2996: data <= 8'h00;
            14'd2997: data <= 8'h00;
            14'd2998: data <= 8'h00;
            14'd2999: data <= 8'h00;
            14'd3000: data <= 8'h00;
            14'd3001: data <= 8'h00;
            14'd3002: data <= 8'h00;
            14'd3003: data <= 8'h00;
            14'd3004: data <= 8'h00;
            14'd3005: data <= 8'h00;
            14'd3006: data <= 8'h0F;
            14'd3007: data <= 8'hFF;
            14'd3008: data <= 8'hFF;
            14'd3009: data <= 8'hFF;
            14'd3010: data <= 8'hFF;
            14'd3011: data <= 8'hFF;
            14'd3012: data <= 8'hFF;
            14'd3013: data <= 8'hFF;
            14'd3014: data <= 8'hFF;
            14'd3015: data <= 8'hFF;
            14'd3016: data <= 8'hFF;
            14'd3017: data <= 8'hFF;
            14'd3018: data <= 8'hFF;
            14'd3019: data <= 8'hFF;
            14'd3020: data <= 8'hFF;
            14'd3021: data <= 8'hFF;
            14'd3022: data <= 8'hFF;
            14'd3023: data <= 8'hFF;
            14'd3024: data <= 8'hFF;
            14'd3025: data <= 8'hFF;
            14'd3026: data <= 8'hFF;
            14'd3027: data <= 8'hFF;
            14'd3028: data <= 8'hFF;
            14'd3029: data <= 8'hFF;
            14'd3030: data <= 8'hFF;
            14'd3031: data <= 8'hFF;
            14'd3032: data <= 8'hFF;
            14'd3033: data <= 8'hF0;
            14'd3034: data <= 8'h00;
            14'd3035: data <= 8'h00;
            14'd3036: data <= 8'h00;
            14'd3037: data <= 8'h00;
            14'd3038: data <= 8'h00;
            14'd3039: data <= 8'h00;
            14'd3040: data <= 8'h00;
            14'd3041: data <= 8'h00;
            14'd3042: data <= 8'h00;
            14'd3043: data <= 8'h00;
            14'd3044: data <= 8'h00;
            14'd3045: data <= 8'h00;
            14'd3046: data <= 8'h0F;
            14'd3047: data <= 8'hFF;
            14'd3048: data <= 8'hFF;
            14'd3049: data <= 8'hFF;
            14'd3050: data <= 8'hFF;
            14'd3051: data <= 8'hFF;
            14'd3052: data <= 8'hFF;
            14'd3053: data <= 8'hFF;
            14'd3054: data <= 8'hFF;
            14'd3055: data <= 8'hFF;
            14'd3056: data <= 8'hFF;
            14'd3057: data <= 8'hFF;
            14'd3058: data <= 8'hFF;
            14'd3059: data <= 8'hFF;
            14'd3060: data <= 8'hFF;
            14'd3061: data <= 8'hFF;
            14'd3062: data <= 8'hFF;
            14'd3063: data <= 8'hFF;
            14'd3064: data <= 8'hFF;
            14'd3065: data <= 8'hFF;
            14'd3066: data <= 8'hFF;
            14'd3067: data <= 8'hFF;
            14'd3068: data <= 8'hFF;
            14'd3069: data <= 8'hFF;
            14'd3070: data <= 8'hFF;
            14'd3071: data <= 8'hFF;
            14'd3072: data <= 8'hFF;
            14'd3073: data <= 8'hF0;
            14'd3074: data <= 8'h00;
            14'd3075: data <= 8'h00;
            14'd3076: data <= 8'h00;
            14'd3077: data <= 8'h00;
            14'd3078: data <= 8'h00;
            14'd3079: data <= 8'h00;
            14'd3080: data <= 8'h00;
            14'd3081: data <= 8'h00;
            14'd3082: data <= 8'h00;
            14'd3083: data <= 8'h00;
            14'd3084: data <= 8'h00;
            14'd3085: data <= 8'h00;
            14'd3086: data <= 8'h0F;
            14'd3087: data <= 8'hFF;
            14'd3088: data <= 8'hFF;
            14'd3089: data <= 8'hFF;
            14'd3090: data <= 8'hFF;
            14'd3091: data <= 8'hFF;
            14'd3092: data <= 8'hFF;
            14'd3093: data <= 8'hFF;
            14'd3094: data <= 8'hFF;
            14'd3095: data <= 8'hFF;
            14'd3096: data <= 8'hFF;
            14'd3097: data <= 8'hFF;
            14'd3098: data <= 8'hFF;
            14'd3099: data <= 8'hFF;
            14'd3100: data <= 8'hFF;
            14'd3101: data <= 8'hFF;
            14'd3102: data <= 8'hFF;
            14'd3103: data <= 8'hFF;
            14'd3104: data <= 8'hFF;
            14'd3105: data <= 8'hFF;
            14'd3106: data <= 8'hFF;
            14'd3107: data <= 8'hFF;
            14'd3108: data <= 8'hFF;
            14'd3109: data <= 8'hFF;
            14'd3110: data <= 8'hFF;
            14'd3111: data <= 8'hFF;
            14'd3112: data <= 8'hFF;
            14'd3113: data <= 8'hF0;
            14'd3114: data <= 8'h00;
            14'd3115: data <= 8'h00;
            14'd3116: data <= 8'h00;
            14'd3117: data <= 8'h00;
            14'd3118: data <= 8'h00;
            14'd3119: data <= 8'h00;
            14'd3120: data <= 8'h00;
            14'd3121: data <= 8'h00;
            14'd3122: data <= 8'h00;
            14'd3123: data <= 8'h00;
            14'd3124: data <= 8'h00;
            14'd3125: data <= 8'h00;
            14'd3126: data <= 8'h0F;
            14'd3127: data <= 8'hFF;
            14'd3128: data <= 8'hFF;
            14'd3129: data <= 8'hFF;
            14'd3130: data <= 8'hFF;
            14'd3131: data <= 8'hFF;
            14'd3132: data <= 8'hFF;
            14'd3133: data <= 8'hFF;
            14'd3134: data <= 8'hFF;
            14'd3135: data <= 8'hFF;
            14'd3136: data <= 8'hFF;
            14'd3137: data <= 8'hE0;
            14'd3138: data <= 8'hFF;
            14'd3139: data <= 8'hFF;
            14'd3140: data <= 8'hFF;
            14'd3141: data <= 8'hFF;
            14'd3142: data <= 8'h83;
            14'd3143: data <= 8'hFF;
            14'd3144: data <= 8'hFF;
            14'd3145: data <= 8'hFF;
            14'd3146: data <= 8'hFF;
            14'd3147: data <= 8'hFF;
            14'd3148: data <= 8'hFF;
            14'd3149: data <= 8'hFF;
            14'd3150: data <= 8'hFF;
            14'd3151: data <= 8'hFF;
            14'd3152: data <= 8'hFF;
            14'd3153: data <= 8'hF0;
            14'd3154: data <= 8'h00;
            14'd3155: data <= 8'h00;
            14'd3156: data <= 8'h00;
            14'd3157: data <= 8'h00;
            14'd3158: data <= 8'h00;
            14'd3159: data <= 8'h00;
            14'd3160: data <= 8'h00;
            14'd3161: data <= 8'h00;
            14'd3162: data <= 8'h00;
            14'd3163: data <= 8'h00;
            14'd3164: data <= 8'h00;
            14'd3165: data <= 8'h00;
            14'd3166: data <= 8'h0F;
            14'd3167: data <= 8'hFF;
            14'd3168: data <= 8'hFF;
            14'd3169: data <= 8'hFF;
            14'd3170: data <= 8'hFF;
            14'd3171: data <= 8'hFF;
            14'd3172: data <= 8'hFF;
            14'd3173: data <= 8'hFF;
            14'd3174: data <= 8'hFF;
            14'd3175: data <= 8'hFF;
            14'd3176: data <= 8'hFF;
            14'd3177: data <= 8'hC0;
            14'd3178: data <= 8'h7F;
            14'd3179: data <= 8'hFF;
            14'd3180: data <= 8'hFF;
            14'd3181: data <= 8'hFF;
            14'd3182: data <= 8'h01;
            14'd3183: data <= 8'hFF;
            14'd3184: data <= 8'hFF;
            14'd3185: data <= 8'hFF;
            14'd3186: data <= 8'hFF;
            14'd3187: data <= 8'hFF;
            14'd3188: data <= 8'hFF;
            14'd3189: data <= 8'hFF;
            14'd3190: data <= 8'hFF;
            14'd3191: data <= 8'hFF;
            14'd3192: data <= 8'hFF;
            14'd3193: data <= 8'hF0;
            14'd3194: data <= 8'h00;
            14'd3195: data <= 8'h00;
            14'd3196: data <= 8'h00;
            14'd3197: data <= 8'h00;
            14'd3198: data <= 8'h00;
            14'd3199: data <= 8'h00;
            14'd3200: data <= 8'h00;
            14'd3201: data <= 8'h00;
            14'd3202: data <= 8'h00;
            14'd3203: data <= 8'h00;
            14'd3204: data <= 8'h00;
            14'd3205: data <= 8'h00;
            14'd3206: data <= 8'h0F;
            14'd3207: data <= 8'hFF;
            14'd3208: data <= 8'hFF;
            14'd3209: data <= 8'hFF;
            14'd3210: data <= 8'hFF;
            14'd3211: data <= 8'hFF;
            14'd3212: data <= 8'hFF;
            14'd3213: data <= 8'hFF;
            14'd3214: data <= 8'hFF;
            14'd3215: data <= 8'hFF;
            14'd3216: data <= 8'hFF;
            14'd3217: data <= 8'h80;
            14'd3218: data <= 8'h3F;
            14'd3219: data <= 8'hFF;
            14'd3220: data <= 8'hFF;
            14'd3221: data <= 8'hFE;
            14'd3222: data <= 8'h01;
            14'd3223: data <= 8'hFF;
            14'd3224: data <= 8'hFF;
            14'd3225: data <= 8'hFF;
            14'd3226: data <= 8'hFF;
            14'd3227: data <= 8'hFF;
            14'd3228: data <= 8'hFF;
            14'd3229: data <= 8'hFF;
            14'd3230: data <= 8'hFF;
            14'd3231: data <= 8'hFF;
            14'd3232: data <= 8'hFF;
            14'd3233: data <= 8'hF0;
            14'd3234: data <= 8'h00;
            14'd3235: data <= 8'h00;
            14'd3236: data <= 8'h00;
            14'd3237: data <= 8'h00;
            14'd3238: data <= 8'h00;
            14'd3239: data <= 8'h00;
            14'd3240: data <= 8'h00;
            14'd3241: data <= 8'h00;
            14'd3242: data <= 8'h00;
            14'd3243: data <= 8'h00;
            14'd3244: data <= 8'h00;
            14'd3245: data <= 8'h00;
            14'd3246: data <= 8'h0F;
            14'd3247: data <= 8'hFF;
            14'd3248: data <= 8'hFF;
            14'd3249: data <= 8'hFF;
            14'd3250: data <= 8'hFF;
            14'd3251: data <= 8'hFF;
            14'd3252: data <= 8'hFF;
            14'd3253: data <= 8'hFF;
            14'd3254: data <= 8'hFF;
            14'd3255: data <= 8'hFF;
            14'd3256: data <= 8'hFF;
            14'd3257: data <= 8'h80;
            14'd3258: data <= 8'h3F;
            14'd3259: data <= 8'hFF;
            14'd3260: data <= 8'hFF;
            14'd3261: data <= 8'hFC;
            14'd3262: data <= 8'h00;
            14'd3263: data <= 8'hFF;
            14'd3264: data <= 8'hFF;
            14'd3265: data <= 8'hFF;
            14'd3266: data <= 8'hFF;
            14'd3267: data <= 8'hFF;
            14'd3268: data <= 8'hFF;
            14'd3269: data <= 8'hFF;
            14'd3270: data <= 8'hFF;
            14'd3271: data <= 8'hFF;
            14'd3272: data <= 8'hFF;
            14'd3273: data <= 8'hF0;
            14'd3274: data <= 8'h00;
            14'd3275: data <= 8'h00;
            14'd3276: data <= 8'h00;
            14'd3277: data <= 8'h00;
            14'd3278: data <= 8'h00;
            14'd3279: data <= 8'h00;
            14'd3280: data <= 8'h00;
            14'd3281: data <= 8'h00;
            14'd3282: data <= 8'h00;
            14'd3283: data <= 8'h00;
            14'd3284: data <= 8'h00;
            14'd3285: data <= 8'h00;
            14'd3286: data <= 8'h0F;
            14'd3287: data <= 8'hFF;
            14'd3288: data <= 8'hFF;
            14'd3289: data <= 8'hFF;
            14'd3290: data <= 8'hFF;
            14'd3291: data <= 8'hFF;
            14'd3292: data <= 8'hFF;
            14'd3293: data <= 8'hFF;
            14'd3294: data <= 8'hFF;
            14'd3295: data <= 8'hFF;
            14'd3296: data <= 8'hFF;
            14'd3297: data <= 8'h00;
            14'd3298: data <= 8'h1F;
            14'd3299: data <= 8'hFF;
            14'd3300: data <= 8'hFF;
            14'd3301: data <= 8'hFC;
            14'd3302: data <= 8'h00;
            14'd3303: data <= 8'hFF;
            14'd3304: data <= 8'hFF;
            14'd3305: data <= 8'hFF;
            14'd3306: data <= 8'hFF;
            14'd3307: data <= 8'hFF;
            14'd3308: data <= 8'hFF;
            14'd3309: data <= 8'hFF;
            14'd3310: data <= 8'hFF;
            14'd3311: data <= 8'hFF;
            14'd3312: data <= 8'hFF;
            14'd3313: data <= 8'hF0;
            14'd3314: data <= 8'h00;
            14'd3315: data <= 8'h00;
            14'd3316: data <= 8'h00;
            14'd3317: data <= 8'h00;
            14'd3318: data <= 8'h00;
            14'd3319: data <= 8'h00;
            14'd3320: data <= 8'h00;
            14'd3321: data <= 8'h00;
            14'd3322: data <= 8'h00;
            14'd3323: data <= 8'h00;
            14'd3324: data <= 8'h00;
            14'd3325: data <= 8'h00;
            14'd3326: data <= 8'h0F;
            14'd3327: data <= 8'hFF;
            14'd3328: data <= 8'hFF;
            14'd3329: data <= 8'hFF;
            14'd3330: data <= 8'hFF;
            14'd3331: data <= 8'hFF;
            14'd3332: data <= 8'hFF;
            14'd3333: data <= 8'hFF;
            14'd3334: data <= 8'hFF;
            14'd3335: data <= 8'hFF;
            14'd3336: data <= 8'hFF;
            14'd3337: data <= 8'h00;
            14'd3338: data <= 8'h1F;
            14'd3339: data <= 8'hFF;
            14'd3340: data <= 8'hFF;
            14'd3341: data <= 8'hF8;
            14'd3342: data <= 8'h00;
            14'd3343: data <= 8'hFF;
            14'd3344: data <= 8'hFF;
            14'd3345: data <= 8'hFF;
            14'd3346: data <= 8'hFF;
            14'd3347: data <= 8'hFF;
            14'd3348: data <= 8'hFF;
            14'd3349: data <= 8'hFF;
            14'd3350: data <= 8'hFF;
            14'd3351: data <= 8'hFF;
            14'd3352: data <= 8'hFF;
            14'd3353: data <= 8'hF0;
            14'd3354: data <= 8'h00;
            14'd3355: data <= 8'h00;
            14'd3356: data <= 8'h00;
            14'd3357: data <= 8'h00;
            14'd3358: data <= 8'h00;
            14'd3359: data <= 8'h00;
            14'd3360: data <= 8'h00;
            14'd3361: data <= 8'h00;
            14'd3362: data <= 8'h00;
            14'd3363: data <= 8'h00;
            14'd3364: data <= 8'h00;
            14'd3365: data <= 8'h00;
            14'd3366: data <= 8'h0F;
            14'd3367: data <= 8'hFF;
            14'd3368: data <= 8'hFF;
            14'd3369: data <= 8'hFF;
            14'd3370: data <= 8'hFF;
            14'd3371: data <= 8'hFF;
            14'd3372: data <= 8'hFF;
            14'd3373: data <= 8'hFF;
            14'd3374: data <= 8'hFF;
            14'd3375: data <= 8'hFF;
            14'd3376: data <= 8'hFF;
            14'd3377: data <= 8'h00;
            14'd3378: data <= 8'h1F;
            14'd3379: data <= 8'hFF;
            14'd3380: data <= 8'hFF;
            14'd3381: data <= 8'hF8;
            14'd3382: data <= 8'h00;
            14'd3383: data <= 8'hFF;
            14'd3384: data <= 8'hFF;
            14'd3385: data <= 8'hFF;
            14'd3386: data <= 8'hFF;
            14'd3387: data <= 8'hFF;
            14'd3388: data <= 8'hFF;
            14'd3389: data <= 8'hFF;
            14'd3390: data <= 8'hFF;
            14'd3391: data <= 8'hFF;
            14'd3392: data <= 8'hFF;
            14'd3393: data <= 8'hF0;
            14'd3394: data <= 8'h00;
            14'd3395: data <= 8'h00;
            14'd3396: data <= 8'h00;
            14'd3397: data <= 8'h00;
            14'd3398: data <= 8'h00;
            14'd3399: data <= 8'h00;
            14'd3400: data <= 8'h00;
            14'd3401: data <= 8'h00;
            14'd3402: data <= 8'h00;
            14'd3403: data <= 8'h00;
            14'd3404: data <= 8'h00;
            14'd3405: data <= 8'h00;
            14'd3406: data <= 8'h0F;
            14'd3407: data <= 8'hFF;
            14'd3408: data <= 8'hFF;
            14'd3409: data <= 8'hFF;
            14'd3410: data <= 8'hFF;
            14'd3411: data <= 8'hFF;
            14'd3412: data <= 8'hFF;
            14'd3413: data <= 8'hFF;
            14'd3414: data <= 8'hFF;
            14'd3415: data <= 8'hFF;
            14'd3416: data <= 8'hFF;
            14'd3417: data <= 8'h00;
            14'd3418: data <= 8'h1F;
            14'd3419: data <= 8'hFF;
            14'd3420: data <= 8'hFF;
            14'd3421: data <= 8'hF8;
            14'd3422: data <= 8'h01;
            14'd3423: data <= 8'hFF;
            14'd3424: data <= 8'hFF;
            14'd3425: data <= 8'hFF;
            14'd3426: data <= 8'hFF;
            14'd3427: data <= 8'hFF;
            14'd3428: data <= 8'hFF;
            14'd3429: data <= 8'hFF;
            14'd3430: data <= 8'hFF;
            14'd3431: data <= 8'hFF;
            14'd3432: data <= 8'hFF;
            14'd3433: data <= 8'hF0;
            14'd3434: data <= 8'h00;
            14'd3435: data <= 8'h00;
            14'd3436: data <= 8'h00;
            14'd3437: data <= 8'h00;
            14'd3438: data <= 8'h00;
            14'd3439: data <= 8'h00;
            14'd3440: data <= 8'h00;
            14'd3441: data <= 8'h00;
            14'd3442: data <= 8'h00;
            14'd3443: data <= 8'h00;
            14'd3444: data <= 8'h00;
            14'd3445: data <= 8'h00;
            14'd3446: data <= 8'h0F;
            14'd3447: data <= 8'hFF;
            14'd3448: data <= 8'hFF;
            14'd3449: data <= 8'hFF;
            14'd3450: data <= 8'hFF;
            14'd3451: data <= 8'hFF;
            14'd3452: data <= 8'hFF;
            14'd3453: data <= 8'hFF;
            14'd3454: data <= 8'hFF;
            14'd3455: data <= 8'hFF;
            14'd3456: data <= 8'hFF;
            14'd3457: data <= 8'h80;
            14'd3458: data <= 8'h3F;
            14'd3459: data <= 8'hFF;
            14'd3460: data <= 8'hFF;
            14'd3461: data <= 8'hFC;
            14'd3462: data <= 8'h01;
            14'd3463: data <= 8'hFF;
            14'd3464: data <= 8'hFF;
            14'd3465: data <= 8'hFF;
            14'd3466: data <= 8'hFF;
            14'd3467: data <= 8'hFF;
            14'd3468: data <= 8'hFF;
            14'd3469: data <= 8'hFF;
            14'd3470: data <= 8'hFF;
            14'd3471: data <= 8'hFF;
            14'd3472: data <= 8'hFF;
            14'd3473: data <= 8'hF0;
            14'd3474: data <= 8'h00;
            14'd3475: data <= 8'h00;
            14'd3476: data <= 8'h00;
            14'd3477: data <= 8'h00;
            14'd3478: data <= 8'h00;
            14'd3479: data <= 8'h00;
            14'd3480: data <= 8'h00;
            14'd3481: data <= 8'h00;
            14'd3482: data <= 8'h00;
            14'd3483: data <= 8'h00;
            14'd3484: data <= 8'h00;
            14'd3485: data <= 8'h00;
            14'd3486: data <= 8'h0F;
            14'd3487: data <= 8'hFF;
            14'd3488: data <= 8'hFF;
            14'd3489: data <= 8'hFF;
            14'd3490: data <= 8'hFF;
            14'd3491: data <= 8'hFF;
            14'd3492: data <= 8'hFF;
            14'd3493: data <= 8'hFF;
            14'd3494: data <= 8'hFF;
            14'd3495: data <= 8'hFF;
            14'd3496: data <= 8'hFF;
            14'd3497: data <= 8'h80;
            14'd3498: data <= 8'h7F;
            14'd3499: data <= 8'hFF;
            14'd3500: data <= 8'hFF;
            14'd3501: data <= 8'hFE;
            14'd3502: data <= 8'h03;
            14'd3503: data <= 8'hFF;
            14'd3504: data <= 8'hFF;
            14'd3505: data <= 8'hFF;
            14'd3506: data <= 8'hFF;
            14'd3507: data <= 8'hFF;
            14'd3508: data <= 8'hFF;
            14'd3509: data <= 8'hFF;
            14'd3510: data <= 8'hFF;
            14'd3511: data <= 8'hFF;
            14'd3512: data <= 8'hFF;
            14'd3513: data <= 8'hF0;
            14'd3514: data <= 8'h00;
            14'd3515: data <= 8'h00;
            14'd3516: data <= 8'h00;
            14'd3517: data <= 8'h00;
            14'd3518: data <= 8'h00;
            14'd3519: data <= 8'h00;
            14'd3520: data <= 8'h00;
            14'd3521: data <= 8'h00;
            14'd3522: data <= 8'h00;
            14'd3523: data <= 8'h00;
            14'd3524: data <= 8'h00;
            14'd3525: data <= 8'h00;
            14'd3526: data <= 8'h0F;
            14'd3527: data <= 8'hFF;
            14'd3528: data <= 8'hFF;
            14'd3529: data <= 8'hFF;
            14'd3530: data <= 8'hFF;
            14'd3531: data <= 8'hFF;
            14'd3532: data <= 8'hFF;
            14'd3533: data <= 8'hFF;
            14'd3534: data <= 8'hFF;
            14'd3535: data <= 8'hFF;
            14'd3536: data <= 8'hFF;
            14'd3537: data <= 8'hC1;
            14'd3538: data <= 8'hFF;
            14'd3539: data <= 8'hFF;
            14'd3540: data <= 8'hFF;
            14'd3541: data <= 8'hFF;
            14'd3542: data <= 8'h0F;
            14'd3543: data <= 8'hFF;
            14'd3544: data <= 8'hFF;
            14'd3545: data <= 8'hFF;
            14'd3546: data <= 8'hFF;
            14'd3547: data <= 8'hFF;
            14'd3548: data <= 8'hFF;
            14'd3549: data <= 8'hFF;
            14'd3550: data <= 8'hFF;
            14'd3551: data <= 8'hFF;
            14'd3552: data <= 8'hFF;
            14'd3553: data <= 8'hF0;
            14'd3554: data <= 8'h00;
            14'd3555: data <= 8'h00;
            14'd3556: data <= 8'h00;
            14'd3557: data <= 8'h00;
            14'd3558: data <= 8'h00;
            14'd3559: data <= 8'h00;
            14'd3560: data <= 8'h00;
            14'd3561: data <= 8'h00;
            14'd3562: data <= 8'h00;
            14'd3563: data <= 8'h00;
            14'd3564: data <= 8'h00;
            14'd3565: data <= 8'h00;
            14'd3566: data <= 8'h0F;
            14'd3567: data <= 8'hFF;
            14'd3568: data <= 8'hFF;
            14'd3569: data <= 8'hFF;
            14'd3570: data <= 8'hFF;
            14'd3571: data <= 8'hFF;
            14'd3572: data <= 8'hFF;
            14'd3573: data <= 8'hFF;
            14'd3574: data <= 8'hFF;
            14'd3575: data <= 8'hFF;
            14'd3576: data <= 8'hFF;
            14'd3577: data <= 8'hF6;
            14'd3578: data <= 8'hFF;
            14'd3579: data <= 8'hFF;
            14'd3580: data <= 8'hFF;
            14'd3581: data <= 8'hFF;
            14'd3582: data <= 8'hFF;
            14'd3583: data <= 8'hFF;
            14'd3584: data <= 8'hFF;
            14'd3585: data <= 8'hFF;
            14'd3586: data <= 8'hFF;
            14'd3587: data <= 8'hFF;
            14'd3588: data <= 8'hFF;
            14'd3589: data <= 8'hFF;
            14'd3590: data <= 8'hFF;
            14'd3591: data <= 8'hFF;
            14'd3592: data <= 8'hFF;
            14'd3593: data <= 8'hF0;
            14'd3594: data <= 8'h00;
            14'd3595: data <= 8'h00;
            14'd3596: data <= 8'h00;
            14'd3597: data <= 8'h00;
            14'd3598: data <= 8'h00;
            14'd3599: data <= 8'h00;
            14'd3600: data <= 8'h00;
            14'd3601: data <= 8'h00;
            14'd3602: data <= 8'h00;
            14'd3603: data <= 8'h00;
            14'd3604: data <= 8'h00;
            14'd3605: data <= 8'h00;
            14'd3606: data <= 8'h0F;
            14'd3607: data <= 8'hFF;
            14'd3608: data <= 8'hFF;
            14'd3609: data <= 8'hFF;
            14'd3610: data <= 8'hFF;
            14'd3611: data <= 8'hFF;
            14'd3612: data <= 8'hFF;
            14'd3613: data <= 8'hFF;
            14'd3614: data <= 8'hFF;
            14'd3615: data <= 8'hFF;
            14'd3616: data <= 8'hFF;
            14'd3617: data <= 8'hFF;
            14'd3618: data <= 8'hFF;
            14'd3619: data <= 8'hFF;
            14'd3620: data <= 8'hFF;
            14'd3621: data <= 8'hFF;
            14'd3622: data <= 8'hFF;
            14'd3623: data <= 8'hFF;
            14'd3624: data <= 8'hFF;
            14'd3625: data <= 8'hFF;
            14'd3626: data <= 8'hFF;
            14'd3627: data <= 8'hFF;
            14'd3628: data <= 8'hFF;
            14'd3629: data <= 8'hFF;
            14'd3630: data <= 8'hFF;
            14'd3631: data <= 8'hFF;
            14'd3632: data <= 8'hFF;
            14'd3633: data <= 8'hF0;
            14'd3634: data <= 8'h00;
            14'd3635: data <= 8'h00;
            14'd3636: data <= 8'h00;
            14'd3637: data <= 8'h00;
            14'd3638: data <= 8'h00;
            14'd3639: data <= 8'h00;
            14'd3640: data <= 8'h00;
            14'd3641: data <= 8'h00;
            14'd3642: data <= 8'h00;
            14'd3643: data <= 8'h00;
            14'd3644: data <= 8'h00;
            14'd3645: data <= 8'h00;
            14'd3646: data <= 8'h0F;
            14'd3647: data <= 8'hFF;
            14'd3648: data <= 8'hFF;
            14'd3649: data <= 8'hFF;
            14'd3650: data <= 8'hFF;
            14'd3651: data <= 8'hFF;
            14'd3652: data <= 8'hFF;
            14'd3653: data <= 8'hFF;
            14'd3654: data <= 8'hFF;
            14'd3655: data <= 8'hFF;
            14'd3656: data <= 8'hFF;
            14'd3657: data <= 8'hFF;
            14'd3658: data <= 8'hFF;
            14'd3659: data <= 8'hFF;
            14'd3660: data <= 8'hFF;
            14'd3661: data <= 8'hFF;
            14'd3662: data <= 8'hFF;
            14'd3663: data <= 8'hFF;
            14'd3664: data <= 8'hFF;
            14'd3665: data <= 8'hFF;
            14'd3666: data <= 8'hFF;
            14'd3667: data <= 8'hFF;
            14'd3668: data <= 8'hFF;
            14'd3669: data <= 8'hFF;
            14'd3670: data <= 8'hFF;
            14'd3671: data <= 8'hFF;
            14'd3672: data <= 8'hFF;
            14'd3673: data <= 8'hF0;
            14'd3674: data <= 8'h00;
            14'd3675: data <= 8'h00;
            14'd3676: data <= 8'h00;
            14'd3677: data <= 8'h00;
            14'd3678: data <= 8'h00;
            14'd3679: data <= 8'h00;
            14'd3680: data <= 8'h00;
            14'd3681: data <= 8'h00;
            14'd3682: data <= 8'h00;
            14'd3683: data <= 8'h00;
            14'd3684: data <= 8'h00;
            14'd3685: data <= 8'h00;
            14'd3686: data <= 8'h0F;
            14'd3687: data <= 8'hFF;
            14'd3688: data <= 8'hFF;
            14'd3689: data <= 8'hFF;
            14'd3690: data <= 8'hFF;
            14'd3691: data <= 8'hFF;
            14'd3692: data <= 8'hFF;
            14'd3693: data <= 8'hFF;
            14'd3694: data <= 8'hFF;
            14'd3695: data <= 8'hFF;
            14'd3696: data <= 8'hFF;
            14'd3697: data <= 8'hFF;
            14'd3698: data <= 8'hFF;
            14'd3699: data <= 8'hFF;
            14'd3700: data <= 8'hFF;
            14'd3701: data <= 8'hFF;
            14'd3702: data <= 8'hFF;
            14'd3703: data <= 8'hFF;
            14'd3704: data <= 8'hFF;
            14'd3705: data <= 8'hFF;
            14'd3706: data <= 8'hFF;
            14'd3707: data <= 8'hFF;
            14'd3708: data <= 8'hFF;
            14'd3709: data <= 8'hFF;
            14'd3710: data <= 8'hFF;
            14'd3711: data <= 8'hFF;
            14'd3712: data <= 8'hFF;
            14'd3713: data <= 8'hF0;
            14'd3714: data <= 8'h00;
            14'd3715: data <= 8'h00;
            14'd3716: data <= 8'h00;
            14'd3717: data <= 8'h00;
            14'd3718: data <= 8'h00;
            14'd3719: data <= 8'h00;
            14'd3720: data <= 8'h00;
            14'd3721: data <= 8'h00;
            14'd3722: data <= 8'h00;
            14'd3723: data <= 8'h00;
            14'd3724: data <= 8'h00;
            14'd3725: data <= 8'h00;
            14'd3726: data <= 8'h0F;
            14'd3727: data <= 8'hFF;
            14'd3728: data <= 8'hFF;
            14'd3729: data <= 8'hFF;
            14'd3730: data <= 8'hFF;
            14'd3731: data <= 8'hFF;
            14'd3732: data <= 8'hFF;
            14'd3733: data <= 8'hFF;
            14'd3734: data <= 8'hFF;
            14'd3735: data <= 8'hFF;
            14'd3736: data <= 8'hFF;
            14'd3737: data <= 8'hFF;
            14'd3738: data <= 8'hFF;
            14'd3739: data <= 8'hFF;
            14'd3740: data <= 8'hFF;
            14'd3741: data <= 8'hFF;
            14'd3742: data <= 8'hFF;
            14'd3743: data <= 8'hFF;
            14'd3744: data <= 8'hFF;
            14'd3745: data <= 8'hFF;
            14'd3746: data <= 8'hFF;
            14'd3747: data <= 8'hFF;
            14'd3748: data <= 8'hFF;
            14'd3749: data <= 8'hFF;
            14'd3750: data <= 8'hFF;
            14'd3751: data <= 8'hFF;
            14'd3752: data <= 8'hFF;
            14'd3753: data <= 8'hF0;
            14'd3754: data <= 8'h00;
            14'd3755: data <= 8'h00;
            14'd3756: data <= 8'h00;
            14'd3757: data <= 8'h00;
            14'd3758: data <= 8'h00;
            14'd3759: data <= 8'h00;
            14'd3760: data <= 8'h00;
            14'd3761: data <= 8'h00;
            14'd3762: data <= 8'h00;
            14'd3763: data <= 8'h00;
            14'd3764: data <= 8'h00;
            14'd3765: data <= 8'h00;
            14'd3766: data <= 8'h0F;
            14'd3767: data <= 8'hFF;
            14'd3768: data <= 8'hFF;
            14'd3769: data <= 8'hFF;
            14'd3770: data <= 8'hFF;
            14'd3771: data <= 8'hFF;
            14'd3772: data <= 8'hFF;
            14'd3773: data <= 8'hFF;
            14'd3774: data <= 8'hFF;
            14'd3775: data <= 8'hFF;
            14'd3776: data <= 8'hFF;
            14'd3777: data <= 8'hFF;
            14'd3778: data <= 8'hFF;
            14'd3779: data <= 8'hFF;
            14'd3780: data <= 8'hFF;
            14'd3781: data <= 8'hFF;
            14'd3782: data <= 8'hFF;
            14'd3783: data <= 8'hFF;
            14'd3784: data <= 8'hFC;
            14'd3785: data <= 8'h7F;
            14'd3786: data <= 8'h8F;
            14'd3787: data <= 8'hFF;
            14'd3788: data <= 8'hFF;
            14'd3789: data <= 8'hFF;
            14'd3790: data <= 8'hFF;
            14'd3791: data <= 8'hFF;
            14'd3792: data <= 8'hFF;
            14'd3793: data <= 8'hF0;
            14'd3794: data <= 8'h00;
            14'd3795: data <= 8'h00;
            14'd3796: data <= 8'h00;
            14'd3797: data <= 8'h00;
            14'd3798: data <= 8'h00;
            14'd3799: data <= 8'h00;
            14'd3800: data <= 8'h00;
            14'd3801: data <= 8'h00;
            14'd3802: data <= 8'h00;
            14'd3803: data <= 8'h00;
            14'd3804: data <= 8'h00;
            14'd3805: data <= 8'h00;
            14'd3806: data <= 8'h0F;
            14'd3807: data <= 8'hFF;
            14'd3808: data <= 8'hFF;
            14'd3809: data <= 8'hFF;
            14'd3810: data <= 8'hFF;
            14'd3811: data <= 8'hFF;
            14'd3812: data <= 8'hFF;
            14'd3813: data <= 8'hFF;
            14'd3814: data <= 8'hFF;
            14'd3815: data <= 8'hFC;
            14'd3816: data <= 8'h3F;
            14'd3817: data <= 8'hFF;
            14'd3818: data <= 8'hFF;
            14'd3819: data <= 8'hFF;
            14'd3820: data <= 8'hFF;
            14'd3821: data <= 8'hFF;
            14'd3822: data <= 8'hFF;
            14'd3823: data <= 8'hFF;
            14'd3824: data <= 8'hF8;
            14'd3825: data <= 8'h3F;
            14'd3826: data <= 8'h0F;
            14'd3827: data <= 8'hFF;
            14'd3828: data <= 8'hFF;
            14'd3829: data <= 8'hFF;
            14'd3830: data <= 8'hFF;
            14'd3831: data <= 8'hFF;
            14'd3832: data <= 8'hFF;
            14'd3833: data <= 8'hF0;
            14'd3834: data <= 8'h00;
            14'd3835: data <= 8'h00;
            14'd3836: data <= 8'h00;
            14'd3837: data <= 8'h00;
            14'd3838: data <= 8'h00;
            14'd3839: data <= 8'h00;
            14'd3840: data <= 8'h00;
            14'd3841: data <= 8'h00;
            14'd3842: data <= 8'h00;
            14'd3843: data <= 8'h00;
            14'd3844: data <= 8'h00;
            14'd3845: data <= 8'h00;
            14'd3846: data <= 8'h0F;
            14'd3847: data <= 8'hFF;
            14'd3848: data <= 8'hFF;
            14'd3849: data <= 8'hFF;
            14'd3850: data <= 8'hFF;
            14'd3851: data <= 8'hFF;
            14'd3852: data <= 8'hFF;
            14'd3853: data <= 8'hFF;
            14'd3854: data <= 8'hFC;
            14'd3855: data <= 8'h3C;
            14'd3856: data <= 8'h1F;
            14'd3857: data <= 8'hFF;
            14'd3858: data <= 8'hFF;
            14'd3859: data <= 8'hFF;
            14'd3860: data <= 8'hFF;
            14'd3861: data <= 8'hFF;
            14'd3862: data <= 8'hFF;
            14'd3863: data <= 8'hFF;
            14'd3864: data <= 8'hF8;
            14'd3865: data <= 8'h3F;
            14'd3866: data <= 8'h0F;
            14'd3867: data <= 8'hFF;
            14'd3868: data <= 8'hFF;
            14'd3869: data <= 8'hFF;
            14'd3870: data <= 8'hFF;
            14'd3871: data <= 8'hFF;
            14'd3872: data <= 8'hFF;
            14'd3873: data <= 8'hF0;
            14'd3874: data <= 8'h00;
            14'd3875: data <= 8'h00;
            14'd3876: data <= 8'h00;
            14'd3877: data <= 8'h00;
            14'd3878: data <= 8'h00;
            14'd3879: data <= 8'h00;
            14'd3880: data <= 8'h00;
            14'd3881: data <= 8'h00;
            14'd3882: data <= 8'h00;
            14'd3883: data <= 8'h00;
            14'd3884: data <= 8'h00;
            14'd3885: data <= 8'h00;
            14'd3886: data <= 8'h0F;
            14'd3887: data <= 8'hFF;
            14'd3888: data <= 8'hFF;
            14'd3889: data <= 8'hFF;
            14'd3890: data <= 8'hFF;
            14'd3891: data <= 8'hFF;
            14'd3892: data <= 8'hFF;
            14'd3893: data <= 8'hFF;
            14'd3894: data <= 8'hF8;
            14'd3895: data <= 8'h18;
            14'd3896: data <= 8'h1F;
            14'd3897: data <= 8'hFF;
            14'd3898: data <= 8'hFF;
            14'd3899: data <= 8'hFF;
            14'd3900: data <= 8'h87;
            14'd3901: data <= 8'hFF;
            14'd3902: data <= 8'hFF;
            14'd3903: data <= 8'hFF;
            14'd3904: data <= 8'hF8;
            14'd3905: data <= 8'h3E;
            14'd3906: data <= 8'h0F;
            14'd3907: data <= 8'hFF;
            14'd3908: data <= 8'hFF;
            14'd3909: data <= 8'hFF;
            14'd3910: data <= 8'hFF;
            14'd3911: data <= 8'hFF;
            14'd3912: data <= 8'hFF;
            14'd3913: data <= 8'hF0;
            14'd3914: data <= 8'h00;
            14'd3915: data <= 8'h00;
            14'd3916: data <= 8'h00;
            14'd3917: data <= 8'h00;
            14'd3918: data <= 8'h00;
            14'd3919: data <= 8'h00;
            14'd3920: data <= 8'h00;
            14'd3921: data <= 8'h00;
            14'd3922: data <= 8'h00;
            14'd3923: data <= 8'h00;
            14'd3924: data <= 8'h00;
            14'd3925: data <= 8'h00;
            14'd3926: data <= 8'h0F;
            14'd3927: data <= 8'hFF;
            14'd3928: data <= 8'hFF;
            14'd3929: data <= 8'hFF;
            14'd3930: data <= 8'hFF;
            14'd3931: data <= 8'hFF;
            14'd3932: data <= 8'hFF;
            14'd3933: data <= 8'hFF;
            14'd3934: data <= 8'hF8;
            14'd3935: data <= 8'h18;
            14'd3936: data <= 8'h0F;
            14'd3937: data <= 8'hFF;
            14'd3938: data <= 8'hFF;
            14'd3939: data <= 8'hFC;
            14'd3940: data <= 8'h00;
            14'd3941: data <= 8'hFF;
            14'd3942: data <= 8'hFF;
            14'd3943: data <= 8'hFF;
            14'd3944: data <= 8'hF8;
            14'd3945: data <= 8'h3E;
            14'd3946: data <= 8'h0F;
            14'd3947: data <= 8'hFF;
            14'd3948: data <= 8'hFF;
            14'd3949: data <= 8'hFF;
            14'd3950: data <= 8'hFF;
            14'd3951: data <= 8'hFF;
            14'd3952: data <= 8'hFF;
            14'd3953: data <= 8'hF0;
            14'd3954: data <= 8'h00;
            14'd3955: data <= 8'h00;
            14'd3956: data <= 8'h00;
            14'd3957: data <= 8'h00;
            14'd3958: data <= 8'h00;
            14'd3959: data <= 8'h00;
            14'd3960: data <= 8'h00;
            14'd3961: data <= 8'h00;
            14'd3962: data <= 8'h00;
            14'd3963: data <= 8'h00;
            14'd3964: data <= 8'h00;
            14'd3965: data <= 8'h00;
            14'd3966: data <= 8'h0F;
            14'd3967: data <= 8'hFF;
            14'd3968: data <= 8'hFF;
            14'd3969: data <= 8'hFF;
            14'd3970: data <= 8'hFF;
            14'd3971: data <= 8'hFF;
            14'd3972: data <= 8'hFF;
            14'd3973: data <= 8'hFF;
            14'd3974: data <= 8'hF8;
            14'd3975: data <= 8'h38;
            14'd3976: data <= 8'h1F;
            14'd3977: data <= 8'hFF;
            14'd3978: data <= 8'hFF;
            14'd3979: data <= 8'hF0;
            14'd3980: data <= 8'h00;
            14'd3981: data <= 8'h7F;
            14'd3982: data <= 8'hFF;
            14'd3983: data <= 8'hFF;
            14'd3984: data <= 8'hF0;
            14'd3985: data <= 8'h3E;
            14'd3986: data <= 8'h0F;
            14'd3987: data <= 8'hFF;
            14'd3988: data <= 8'hFF;
            14'd3989: data <= 8'hFF;
            14'd3990: data <= 8'hFF;
            14'd3991: data <= 8'hFF;
            14'd3992: data <= 8'hFF;
            14'd3993: data <= 8'hF0;
            14'd3994: data <= 8'h00;
            14'd3995: data <= 8'h00;
            14'd3996: data <= 8'h00;
            14'd3997: data <= 8'h00;
            14'd3998: data <= 8'h00;
            14'd3999: data <= 8'h00;
            14'd4000: data <= 8'h00;
            14'd4001: data <= 8'h00;
            14'd4002: data <= 8'h00;
            14'd4003: data <= 8'h00;
            14'd4004: data <= 8'h00;
            14'd4005: data <= 8'h00;
            14'd4006: data <= 8'h0F;
            14'd4007: data <= 8'hFF;
            14'd4008: data <= 8'hF7;
            14'd4009: data <= 8'hFF;
            14'd4010: data <= 8'hFF;
            14'd4011: data <= 8'hFF;
            14'd4012: data <= 8'hFF;
            14'd4013: data <= 8'hFF;
            14'd4014: data <= 8'hF0;
            14'd4015: data <= 8'h38;
            14'd4016: data <= 8'h1F;
            14'd4017: data <= 8'hFF;
            14'd4018: data <= 8'hFF;
            14'd4019: data <= 8'hE0;
            14'd4020: data <= 8'h00;
            14'd4021: data <= 8'h3F;
            14'd4022: data <= 8'hFF;
            14'd4023: data <= 8'hFF;
            14'd4024: data <= 8'hF8;
            14'd4025: data <= 8'h7E;
            14'd4026: data <= 8'h0F;
            14'd4027: data <= 8'hFF;
            14'd4028: data <= 8'hFF;
            14'd4029: data <= 8'hFF;
            14'd4030: data <= 8'hFF;
            14'd4031: data <= 8'hFF;
            14'd4032: data <= 8'hFF;
            14'd4033: data <= 8'hF0;
            14'd4034: data <= 8'h00;
            14'd4035: data <= 8'h00;
            14'd4036: data <= 8'h00;
            14'd4037: data <= 8'h00;
            14'd4038: data <= 8'h00;
            14'd4039: data <= 8'h00;
            14'd4040: data <= 8'h00;
            14'd4041: data <= 8'h00;
            14'd4042: data <= 8'h00;
            14'd4043: data <= 8'h00;
            14'd4044: data <= 8'h00;
            14'd4045: data <= 8'h00;
            14'd4046: data <= 8'h0F;
            14'd4047: data <= 8'hFF;
            14'd4048: data <= 8'hFF;
            14'd4049: data <= 8'hFF;
            14'd4050: data <= 8'hFF;
            14'd4051: data <= 8'hFF;
            14'd4052: data <= 8'hFF;
            14'd4053: data <= 8'hFF;
            14'd4054: data <= 8'hF8;
            14'd4055: data <= 8'h38;
            14'd4056: data <= 8'h3F;
            14'd4057: data <= 8'hFF;
            14'd4058: data <= 8'hFF;
            14'd4059: data <= 8'hC0;
            14'd4060: data <= 8'h00;
            14'd4061: data <= 8'h1F;
            14'd4062: data <= 8'hFF;
            14'd4063: data <= 8'hFF;
            14'd4064: data <= 8'hF8;
            14'd4065: data <= 8'hFF;
            14'd4066: data <= 8'h1F;
            14'd4067: data <= 8'hFF;
            14'd4068: data <= 8'hFF;
            14'd4069: data <= 8'hFF;
            14'd4070: data <= 8'hFF;
            14'd4071: data <= 8'hFF;
            14'd4072: data <= 8'hFF;
            14'd4073: data <= 8'hF0;
            14'd4074: data <= 8'h00;
            14'd4075: data <= 8'h00;
            14'd4076: data <= 8'h00;
            14'd4077: data <= 8'h00;
            14'd4078: data <= 8'h00;
            14'd4079: data <= 8'h00;
            14'd4080: data <= 8'h00;
            14'd4081: data <= 8'h00;
            14'd4082: data <= 8'h00;
            14'd4083: data <= 8'h00;
            14'd4084: data <= 8'h00;
            14'd4085: data <= 8'h00;
            14'd4086: data <= 8'h0F;
            14'd4087: data <= 8'hFF;
            14'd4088: data <= 8'hFF;
            14'd4089: data <= 8'hFF;
            14'd4090: data <= 8'hFF;
            14'd4091: data <= 8'hFF;
            14'd4092: data <= 8'hFF;
            14'd4093: data <= 8'hFF;
            14'd4094: data <= 8'hF8;
            14'd4095: data <= 8'h78;
            14'd4096: data <= 8'h3F;
            14'd4097: data <= 8'hFF;
            14'd4098: data <= 8'hFF;
            14'd4099: data <= 8'h00;
            14'd4100: data <= 8'h00;
            14'd4101: data <= 8'h0F;
            14'd4102: data <= 8'hFF;
            14'd4103: data <= 8'hFC;
            14'd4104: data <= 8'hFD;
            14'd4105: data <= 8'hFF;
            14'd4106: data <= 8'hFF;
            14'd4107: data <= 8'hFF;
            14'd4108: data <= 8'hFF;
            14'd4109: data <= 8'hFF;
            14'd4110: data <= 8'hFF;
            14'd4111: data <= 8'hFF;
            14'd4112: data <= 8'hFF;
            14'd4113: data <= 8'hF0;
            14'd4114: data <= 8'h00;
            14'd4115: data <= 8'h00;
            14'd4116: data <= 8'h00;
            14'd4117: data <= 8'h00;
            14'd4118: data <= 8'h00;
            14'd4119: data <= 8'h00;
            14'd4120: data <= 8'h00;
            14'd4121: data <= 8'h00;
            14'd4122: data <= 8'h00;
            14'd4123: data <= 8'h00;
            14'd4124: data <= 8'h00;
            14'd4125: data <= 8'h00;
            14'd4126: data <= 8'h0F;
            14'd4127: data <= 8'hFF;
            14'd4128: data <= 8'hFF;
            14'd4129: data <= 8'hFF;
            14'd4130: data <= 8'hFF;
            14'd4131: data <= 8'hFF;
            14'd4132: data <= 8'hFF;
            14'd4133: data <= 8'hFF;
            14'd4134: data <= 8'hF8;
            14'd4135: data <= 8'h78;
            14'd4136: data <= 8'hFF;
            14'd4137: data <= 8'hFF;
            14'd4138: data <= 8'hFE;
            14'd4139: data <= 8'h00;
            14'd4140: data <= 8'h60;
            14'd4141: data <= 8'h03;
            14'd4142: data <= 8'hFF;
            14'd4143: data <= 8'hF0;
            14'd4144: data <= 8'h7F;
            14'd4145: data <= 8'hFF;
            14'd4146: data <= 8'hFF;
            14'd4147: data <= 8'hFF;
            14'd4148: data <= 8'hFF;
            14'd4149: data <= 8'hFF;
            14'd4150: data <= 8'hFF;
            14'd4151: data <= 8'hFF;
            14'd4152: data <= 8'hFF;
            14'd4153: data <= 8'hF0;
            14'd4154: data <= 8'h00;
            14'd4155: data <= 8'h00;
            14'd4156: data <= 8'h00;
            14'd4157: data <= 8'h00;
            14'd4158: data <= 8'h00;
            14'd4159: data <= 8'h00;
            14'd4160: data <= 8'h00;
            14'd4161: data <= 8'h00;
            14'd4162: data <= 8'h00;
            14'd4163: data <= 8'h00;
            14'd4164: data <= 8'h00;
            14'd4165: data <= 8'h00;
            14'd4166: data <= 8'h0F;
            14'd4167: data <= 8'hFF;
            14'd4168: data <= 8'hFF;
            14'd4169: data <= 8'hFF;
            14'd4170: data <= 8'hFF;
            14'd4171: data <= 8'hFF;
            14'd4172: data <= 8'hFF;
            14'd4173: data <= 8'hFF;
            14'd4174: data <= 8'hFC;
            14'd4175: data <= 8'hFF;
            14'd4176: data <= 8'hFF;
            14'd4177: data <= 8'hFF;
            14'd4178: data <= 8'hFE;
            14'd4179: data <= 8'h01;
            14'd4180: data <= 8'hF8;
            14'd4181: data <= 8'h03;
            14'd4182: data <= 8'hFF;
            14'd4183: data <= 8'hF0;
            14'd4184: data <= 8'h7F;
            14'd4185: data <= 8'hFF;
            14'd4186: data <= 8'hFF;
            14'd4187: data <= 8'hFF;
            14'd4188: data <= 8'hFF;
            14'd4189: data <= 8'hFF;
            14'd4190: data <= 8'hFF;
            14'd4191: data <= 8'hFF;
            14'd4192: data <= 8'hFF;
            14'd4193: data <= 8'hF0;
            14'd4194: data <= 8'h00;
            14'd4195: data <= 8'h00;
            14'd4196: data <= 8'h00;
            14'd4197: data <= 8'h00;
            14'd4198: data <= 8'h00;
            14'd4199: data <= 8'h00;
            14'd4200: data <= 8'h00;
            14'd4201: data <= 8'h00;
            14'd4202: data <= 8'h00;
            14'd4203: data <= 8'h00;
            14'd4204: data <= 8'h00;
            14'd4205: data <= 8'h00;
            14'd4206: data <= 8'h0F;
            14'd4207: data <= 8'hFF;
            14'd4208: data <= 8'hFF;
            14'd4209: data <= 8'hFF;
            14'd4210: data <= 8'hFF;
            14'd4211: data <= 8'hFF;
            14'd4212: data <= 8'hFF;
            14'd4213: data <= 8'hFF;
            14'd4214: data <= 8'hFF;
            14'd4215: data <= 8'hFF;
            14'd4216: data <= 8'hFF;
            14'd4217: data <= 8'hFF;
            14'd4218: data <= 8'hFC;
            14'd4219: data <= 8'h07;
            14'd4220: data <= 8'hFE;
            14'd4221: data <= 8'h03;
            14'd4222: data <= 8'hFF;
            14'd4223: data <= 8'hE0;
            14'd4224: data <= 8'h7F;
            14'd4225: data <= 8'hFF;
            14'd4226: data <= 8'hFF;
            14'd4227: data <= 8'hFF;
            14'd4228: data <= 8'hFF;
            14'd4229: data <= 8'hFF;
            14'd4230: data <= 8'hFF;
            14'd4231: data <= 8'hFF;
            14'd4232: data <= 8'hFF;
            14'd4233: data <= 8'hF0;
            14'd4234: data <= 8'h00;
            14'd4235: data <= 8'h00;
            14'd4236: data <= 8'h00;
            14'd4237: data <= 8'h00;
            14'd4238: data <= 8'h00;
            14'd4239: data <= 8'h00;
            14'd4240: data <= 8'h00;
            14'd4241: data <= 8'h00;
            14'd4242: data <= 8'h00;
            14'd4243: data <= 8'h00;
            14'd4244: data <= 8'h00;
            14'd4245: data <= 8'h00;
            14'd4246: data <= 8'h0F;
            14'd4247: data <= 8'hFF;
            14'd4248: data <= 8'hFF;
            14'd4249: data <= 8'hFF;
            14'd4250: data <= 8'hFF;
            14'd4251: data <= 8'hFF;
            14'd4252: data <= 8'hFF;
            14'd4253: data <= 8'hFF;
            14'd4254: data <= 8'hFF;
            14'd4255: data <= 8'hFF;
            14'd4256: data <= 8'hFF;
            14'd4257: data <= 8'hFF;
            14'd4258: data <= 8'hFC;
            14'd4259: data <= 8'h0F;
            14'd4260: data <= 8'hFF;
            14'd4261: data <= 8'h01;
            14'd4262: data <= 8'hFF;
            14'd4263: data <= 8'hC0;
            14'd4264: data <= 8'h7F;
            14'd4265: data <= 8'hFF;
            14'd4266: data <= 8'hFF;
            14'd4267: data <= 8'hFF;
            14'd4268: data <= 8'hFF;
            14'd4269: data <= 8'hFF;
            14'd4270: data <= 8'hFF;
            14'd4271: data <= 8'hFF;
            14'd4272: data <= 8'hFF;
            14'd4273: data <= 8'hF0;
            14'd4274: data <= 8'h00;
            14'd4275: data <= 8'h00;
            14'd4276: data <= 8'h00;
            14'd4277: data <= 8'h00;
            14'd4278: data <= 8'h00;
            14'd4279: data <= 8'h00;
            14'd4280: data <= 8'h00;
            14'd4281: data <= 8'h00;
            14'd4282: data <= 8'h00;
            14'd4283: data <= 8'h00;
            14'd4284: data <= 8'h00;
            14'd4285: data <= 8'h00;
            14'd4286: data <= 8'h0F;
            14'd4287: data <= 8'hFF;
            14'd4288: data <= 8'hFF;
            14'd4289: data <= 8'hFF;
            14'd4290: data <= 8'hFF;
            14'd4291: data <= 8'hFF;
            14'd4292: data <= 8'hFF;
            14'd4293: data <= 8'hFF;
            14'd4294: data <= 8'hFF;
            14'd4295: data <= 8'hFF;
            14'd4296: data <= 8'hFF;
            14'd4297: data <= 8'hFF;
            14'd4298: data <= 8'hFC;
            14'd4299: data <= 8'h1F;
            14'd4300: data <= 8'hFF;
            14'd4301: data <= 8'h83;
            14'd4302: data <= 8'hFF;
            14'd4303: data <= 8'hC0;
            14'd4304: data <= 8'hFF;
            14'd4305: data <= 8'hFF;
            14'd4306: data <= 8'hFF;
            14'd4307: data <= 8'hFF;
            14'd4308: data <= 8'hFF;
            14'd4309: data <= 8'hFF;
            14'd4310: data <= 8'hFF;
            14'd4311: data <= 8'hFF;
            14'd4312: data <= 8'hFF;
            14'd4313: data <= 8'hF0;
            14'd4314: data <= 8'h00;
            14'd4315: data <= 8'h00;
            14'd4316: data <= 8'h00;
            14'd4317: data <= 8'h00;
            14'd4318: data <= 8'h00;
            14'd4319: data <= 8'h00;
            14'd4320: data <= 8'h00;
            14'd4321: data <= 8'h00;
            14'd4322: data <= 8'h00;
            14'd4323: data <= 8'h00;
            14'd4324: data <= 8'h00;
            14'd4325: data <= 8'h00;
            14'd4326: data <= 8'h0F;
            14'd4327: data <= 8'hFF;
            14'd4328: data <= 8'hFF;
            14'd4329: data <= 8'hFF;
            14'd4330: data <= 8'hFF;
            14'd4331: data <= 8'hFF;
            14'd4332: data <= 8'hFF;
            14'd4333: data <= 8'hFF;
            14'd4334: data <= 8'hFF;
            14'd4335: data <= 8'hFF;
            14'd4336: data <= 8'hFF;
            14'd4337: data <= 8'hFF;
            14'd4338: data <= 8'hF8;
            14'd4339: data <= 8'h3F;
            14'd4340: data <= 8'hFF;
            14'd4341: data <= 8'hE7;
            14'd4342: data <= 8'hFF;
            14'd4343: data <= 8'h81;
            14'd4344: data <= 8'hFF;
            14'd4345: data <= 8'hFF;
            14'd4346: data <= 8'hFF;
            14'd4347: data <= 8'hFF;
            14'd4348: data <= 8'hFF;
            14'd4349: data <= 8'hFF;
            14'd4350: data <= 8'hFF;
            14'd4351: data <= 8'hFF;
            14'd4352: data <= 8'hFF;
            14'd4353: data <= 8'hF0;
            14'd4354: data <= 8'h00;
            14'd4355: data <= 8'h00;
            14'd4356: data <= 8'h00;
            14'd4357: data <= 8'h00;
            14'd4358: data <= 8'h00;
            14'd4359: data <= 8'h00;
            14'd4360: data <= 8'h00;
            14'd4361: data <= 8'h00;
            14'd4362: data <= 8'h00;
            14'd4363: data <= 8'h00;
            14'd4364: data <= 8'h00;
            14'd4365: data <= 8'h00;
            14'd4366: data <= 8'h0F;
            14'd4367: data <= 8'hFF;
            14'd4368: data <= 8'hFF;
            14'd4369: data <= 8'hFF;
            14'd4370: data <= 8'hFF;
            14'd4371: data <= 8'hFF;
            14'd4372: data <= 8'hFF;
            14'd4373: data <= 8'hFF;
            14'd4374: data <= 8'hFF;
            14'd4375: data <= 8'hFF;
            14'd4376: data <= 8'hFF;
            14'd4377: data <= 8'hFF;
            14'd4378: data <= 8'hF8;
            14'd4379: data <= 8'h3F;
            14'd4380: data <= 8'hFF;
            14'd4381: data <= 8'hFF;
            14'd4382: data <= 8'hFF;
            14'd4383: data <= 8'h81;
            14'd4384: data <= 8'hFF;
            14'd4385: data <= 8'hFF;
            14'd4386: data <= 8'hFF;
            14'd4387: data <= 8'hFF;
            14'd4388: data <= 8'hFF;
            14'd4389: data <= 8'hFF;
            14'd4390: data <= 8'hFF;
            14'd4391: data <= 8'hFF;
            14'd4392: data <= 8'hFF;
            14'd4393: data <= 8'hF0;
            14'd4394: data <= 8'h00;
            14'd4395: data <= 8'h00;
            14'd4396: data <= 8'h00;
            14'd4397: data <= 8'h00;
            14'd4398: data <= 8'h00;
            14'd4399: data <= 8'h00;
            14'd4400: data <= 8'h00;
            14'd4401: data <= 8'h00;
            14'd4402: data <= 8'h00;
            14'd4403: data <= 8'h00;
            14'd4404: data <= 8'h00;
            14'd4405: data <= 8'h00;
            14'd4406: data <= 8'h0F;
            14'd4407: data <= 8'hEF;
            14'd4408: data <= 8'hFF;
            14'd4409: data <= 8'hFF;
            14'd4410: data <= 8'hFF;
            14'd4411: data <= 8'hFF;
            14'd4412: data <= 8'hFF;
            14'd4413: data <= 8'hFF;
            14'd4414: data <= 8'hFF;
            14'd4415: data <= 8'hFF;
            14'd4416: data <= 8'hFF;
            14'd4417: data <= 8'hFF;
            14'd4418: data <= 8'hFE;
            14'd4419: data <= 8'hFF;
            14'd4420: data <= 8'hFF;
            14'd4421: data <= 8'hFF;
            14'd4422: data <= 8'hFF;
            14'd4423: data <= 8'h03;
            14'd4424: data <= 8'hFF;
            14'd4425: data <= 8'hFF;
            14'd4426: data <= 8'hFF;
            14'd4427: data <= 8'hFF;
            14'd4428: data <= 8'hFF;
            14'd4429: data <= 8'hFF;
            14'd4430: data <= 8'hFF;
            14'd4431: data <= 8'hFF;
            14'd4432: data <= 8'hFF;
            14'd4433: data <= 8'hF0;
            14'd4434: data <= 8'h00;
            14'd4435: data <= 8'h00;
            14'd4436: data <= 8'h00;
            14'd4437: data <= 8'h00;
            14'd4438: data <= 8'h00;
            14'd4439: data <= 8'h00;
            14'd4440: data <= 8'h00;
            14'd4441: data <= 8'h00;
            14'd4442: data <= 8'h00;
            14'd4443: data <= 8'h00;
            14'd4444: data <= 8'h00;
            14'd4445: data <= 8'h00;
            14'd4446: data <= 8'h0F;
            14'd4447: data <= 8'hFF;
            14'd4448: data <= 8'hFF;
            14'd4449: data <= 8'hFF;
            14'd4450: data <= 8'hFF;
            14'd4451: data <= 8'hFF;
            14'd4452: data <= 8'hFF;
            14'd4453: data <= 8'hFF;
            14'd4454: data <= 8'hFF;
            14'd4455: data <= 8'hFF;
            14'd4456: data <= 8'hFF;
            14'd4457: data <= 8'hFF;
            14'd4458: data <= 8'hFF;
            14'd4459: data <= 8'hFF;
            14'd4460: data <= 8'hFF;
            14'd4461: data <= 8'hFF;
            14'd4462: data <= 8'hFE;
            14'd4463: data <= 8'h03;
            14'd4464: data <= 8'hFF;
            14'd4465: data <= 8'hFF;
            14'd4466: data <= 8'hFF;
            14'd4467: data <= 8'hFF;
            14'd4468: data <= 8'hFF;
            14'd4469: data <= 8'hFF;
            14'd4470: data <= 8'hFF;
            14'd4471: data <= 8'hFF;
            14'd4472: data <= 8'hFF;
            14'd4473: data <= 8'hF0;
            14'd4474: data <= 8'h00;
            14'd4475: data <= 8'h00;
            14'd4476: data <= 8'h00;
            14'd4477: data <= 8'h00;
            14'd4478: data <= 8'h00;
            14'd4479: data <= 8'h00;
            14'd4480: data <= 8'h00;
            14'd4481: data <= 8'h00;
            14'd4482: data <= 8'h00;
            14'd4483: data <= 8'h00;
            14'd4484: data <= 8'h00;
            14'd4485: data <= 8'h00;
            14'd4486: data <= 8'h0F;
            14'd4487: data <= 8'hFF;
            14'd4488: data <= 8'hFF;
            14'd4489: data <= 8'hFF;
            14'd4490: data <= 8'hFF;
            14'd4491: data <= 8'hFF;
            14'd4492: data <= 8'hFF;
            14'd4493: data <= 8'hFF;
            14'd4494: data <= 8'hFF;
            14'd4495: data <= 8'hFF;
            14'd4496: data <= 8'hFF;
            14'd4497: data <= 8'hFF;
            14'd4498: data <= 8'hFF;
            14'd4499: data <= 8'hFF;
            14'd4500: data <= 8'hFF;
            14'd4501: data <= 8'hFF;
            14'd4502: data <= 8'hFE;
            14'd4503: data <= 8'h07;
            14'd4504: data <= 8'hFF;
            14'd4505: data <= 8'hFF;
            14'd4506: data <= 8'hFF;
            14'd4507: data <= 8'hFF;
            14'd4508: data <= 8'hFF;
            14'd4509: data <= 8'hFF;
            14'd4510: data <= 8'hFF;
            14'd4511: data <= 8'hFF;
            14'd4512: data <= 8'hFF;
            14'd4513: data <= 8'hF0;
            14'd4514: data <= 8'h00;
            14'd4515: data <= 8'h00;
            14'd4516: data <= 8'h00;
            14'd4517: data <= 8'h00;
            14'd4518: data <= 8'h00;
            14'd4519: data <= 8'h00;
            14'd4520: data <= 8'h00;
            14'd4521: data <= 8'h00;
            14'd4522: data <= 8'h00;
            14'd4523: data <= 8'h00;
            14'd4524: data <= 8'h00;
            14'd4525: data <= 8'h00;
            14'd4526: data <= 8'h0F;
            14'd4527: data <= 8'hFF;
            14'd4528: data <= 8'hFF;
            14'd4529: data <= 8'hFF;
            14'd4530: data <= 8'hFF;
            14'd4531: data <= 8'hFF;
            14'd4532: data <= 8'hFF;
            14'd4533: data <= 8'hFF;
            14'd4534: data <= 8'hFF;
            14'd4535: data <= 8'hFF;
            14'd4536: data <= 8'hFF;
            14'd4537: data <= 8'hFF;
            14'd4538: data <= 8'hFF;
            14'd4539: data <= 8'hFF;
            14'd4540: data <= 8'hFF;
            14'd4541: data <= 8'hFF;
            14'd4542: data <= 8'hFE;
            14'd4543: data <= 8'h0F;
            14'd4544: data <= 8'hFF;
            14'd4545: data <= 8'hE1;
            14'd4546: data <= 8'hFF;
            14'd4547: data <= 8'hFF;
            14'd4548: data <= 8'hFF;
            14'd4549: data <= 8'hFF;
            14'd4550: data <= 8'hFF;
            14'd4551: data <= 8'hFF;
            14'd4552: data <= 8'hFF;
            14'd4553: data <= 8'hF0;
            14'd4554: data <= 8'h00;
            14'd4555: data <= 8'h00;
            14'd4556: data <= 8'h00;
            14'd4557: data <= 8'h00;
            14'd4558: data <= 8'h00;
            14'd4559: data <= 8'h00;
            14'd4560: data <= 8'h00;
            14'd4561: data <= 8'h00;
            14'd4562: data <= 8'h00;
            14'd4563: data <= 8'h00;
            14'd4564: data <= 8'h00;
            14'd4565: data <= 8'h00;
            14'd4566: data <= 8'h0F;
            14'd4567: data <= 8'hFF;
            14'd4568: data <= 8'hFF;
            14'd4569: data <= 8'hFF;
            14'd4570: data <= 8'hFF;
            14'd4571: data <= 8'hFF;
            14'd4572: data <= 8'hFF;
            14'd4573: data <= 8'hFF;
            14'd4574: data <= 8'hFF;
            14'd4575: data <= 8'hFF;
            14'd4576: data <= 8'hFF;
            14'd4577: data <= 8'hFF;
            14'd4578: data <= 8'hFF;
            14'd4579: data <= 8'hFF;
            14'd4580: data <= 8'hFF;
            14'd4581: data <= 8'hFF;
            14'd4582: data <= 8'hFC;
            14'd4583: data <= 8'h0F;
            14'd4584: data <= 8'hFF;
            14'd4585: data <= 8'hC1;
            14'd4586: data <= 8'hFF;
            14'd4587: data <= 8'hFF;
            14'd4588: data <= 8'hFF;
            14'd4589: data <= 8'hFF;
            14'd4590: data <= 8'hFF;
            14'd4591: data <= 8'hFF;
            14'd4592: data <= 8'hFF;
            14'd4593: data <= 8'hF0;
            14'd4594: data <= 8'h00;
            14'd4595: data <= 8'h00;
            14'd4596: data <= 8'h00;
            14'd4597: data <= 8'h00;
            14'd4598: data <= 8'h00;
            14'd4599: data <= 8'h00;
            14'd4600: data <= 8'h00;
            14'd4601: data <= 8'h00;
            14'd4602: data <= 8'h00;
            14'd4603: data <= 8'h00;
            14'd4604: data <= 8'h00;
            14'd4605: data <= 8'h00;
            14'd4606: data <= 8'h0F;
            14'd4607: data <= 8'hFF;
            14'd4608: data <= 8'hFF;
            14'd4609: data <= 8'hFF;
            14'd4610: data <= 8'hFF;
            14'd4611: data <= 8'hFF;
            14'd4612: data <= 8'hFF;
            14'd4613: data <= 8'hFF;
            14'd4614: data <= 8'hFF;
            14'd4615: data <= 8'hFF;
            14'd4616: data <= 8'hFF;
            14'd4617: data <= 8'hFF;
            14'd4618: data <= 8'hFF;
            14'd4619: data <= 8'hFF;
            14'd4620: data <= 8'hFF;
            14'd4621: data <= 8'hFF;
            14'd4622: data <= 8'hF8;
            14'd4623: data <= 8'h0F;
            14'd4624: data <= 8'hFF;
            14'd4625: data <= 8'h81;
            14'd4626: data <= 8'hFF;
            14'd4627: data <= 8'hFF;
            14'd4628: data <= 8'hFF;
            14'd4629: data <= 8'hFF;
            14'd4630: data <= 8'hFF;
            14'd4631: data <= 8'hFF;
            14'd4632: data <= 8'hFF;
            14'd4633: data <= 8'hF0;
            14'd4634: data <= 8'h00;
            14'd4635: data <= 8'h00;
            14'd4636: data <= 8'h00;
            14'd4637: data <= 8'h00;
            14'd4638: data <= 8'h00;
            14'd4639: data <= 8'h00;
            14'd4640: data <= 8'h00;
            14'd4641: data <= 8'h00;
            14'd4642: data <= 8'h00;
            14'd4643: data <= 8'h00;
            14'd4644: data <= 8'h00;
            14'd4645: data <= 8'h00;
            14'd4646: data <= 8'h0F;
            14'd4647: data <= 8'hFF;
            14'd4648: data <= 8'hFF;
            14'd4649: data <= 8'hFF;
            14'd4650: data <= 8'hFF;
            14'd4651: data <= 8'hFF;
            14'd4652: data <= 8'hFF;
            14'd4653: data <= 8'hFF;
            14'd4654: data <= 8'hFF;
            14'd4655: data <= 8'hFF;
            14'd4656: data <= 8'hFF;
            14'd4657: data <= 8'hFF;
            14'd4658: data <= 8'hFF;
            14'd4659: data <= 8'hFE;
            14'd4660: data <= 8'hFF;
            14'd4661: data <= 8'hFF;
            14'd4662: data <= 8'hF8;
            14'd4663: data <= 8'h1F;
            14'd4664: data <= 8'hFF;
            14'd4665: data <= 8'h03;
            14'd4666: data <= 8'hFF;
            14'd4667: data <= 8'hFF;
            14'd4668: data <= 8'hFF;
            14'd4669: data <= 8'hFF;
            14'd4670: data <= 8'hFF;
            14'd4671: data <= 8'hFF;
            14'd4672: data <= 8'hFF;
            14'd4673: data <= 8'hF0;
            14'd4674: data <= 8'h00;
            14'd4675: data <= 8'h00;
            14'd4676: data <= 8'h00;
            14'd4677: data <= 8'h00;
            14'd4678: data <= 8'h00;
            14'd4679: data <= 8'h00;
            14'd4680: data <= 8'h00;
            14'd4681: data <= 8'h00;
            14'd4682: data <= 8'h00;
            14'd4683: data <= 8'h00;
            14'd4684: data <= 8'h00;
            14'd4685: data <= 8'h00;
            14'd4686: data <= 8'h0F;
            14'd4687: data <= 8'hFF;
            14'd4688: data <= 8'hFF;
            14'd4689: data <= 8'hFF;
            14'd4690: data <= 8'hFF;
            14'd4691: data <= 8'hFF;
            14'd4692: data <= 8'hFF;
            14'd4693: data <= 8'hFF;
            14'd4694: data <= 8'hFF;
            14'd4695: data <= 8'hFF;
            14'd4696: data <= 8'hFF;
            14'd4697: data <= 8'hFF;
            14'd4698: data <= 8'hFF;
            14'd4699: data <= 8'hFF;
            14'd4700: data <= 8'hFF;
            14'd4701: data <= 8'hFF;
            14'd4702: data <= 8'hF0;
            14'd4703: data <= 8'h1F;
            14'd4704: data <= 8'hFE;
            14'd4705: data <= 8'h03;
            14'd4706: data <= 8'hFF;
            14'd4707: data <= 8'hFF;
            14'd4708: data <= 8'hFF;
            14'd4709: data <= 8'hFF;
            14'd4710: data <= 8'hFF;
            14'd4711: data <= 8'hFF;
            14'd4712: data <= 8'hFF;
            14'd4713: data <= 8'hF0;
            14'd4714: data <= 8'h00;
            14'd4715: data <= 8'h00;
            14'd4716: data <= 8'h00;
            14'd4717: data <= 8'h00;
            14'd4718: data <= 8'h00;
            14'd4719: data <= 8'h00;
            14'd4720: data <= 8'h00;
            14'd4721: data <= 8'h00;
            14'd4722: data <= 8'h00;
            14'd4723: data <= 8'h00;
            14'd4724: data <= 8'h00;
            14'd4725: data <= 8'h00;
            14'd4726: data <= 8'h0F;
            14'd4727: data <= 8'hFF;
            14'd4728: data <= 8'hFF;
            14'd4729: data <= 8'hFF;
            14'd4730: data <= 8'hFF;
            14'd4731: data <= 8'hFF;
            14'd4732: data <= 8'hFF;
            14'd4733: data <= 8'hFF;
            14'd4734: data <= 8'hFF;
            14'd4735: data <= 8'hFF;
            14'd4736: data <= 8'hFF;
            14'd4737: data <= 8'hFF;
            14'd4738: data <= 8'hFF;
            14'd4739: data <= 8'hFF;
            14'd4740: data <= 8'hFF;
            14'd4741: data <= 8'hFF;
            14'd4742: data <= 8'hF0;
            14'd4743: data <= 8'h3F;
            14'd4744: data <= 8'hFE;
            14'd4745: data <= 8'h07;
            14'd4746: data <= 8'hFF;
            14'd4747: data <= 8'hFF;
            14'd4748: data <= 8'hFF;
            14'd4749: data <= 8'hFF;
            14'd4750: data <= 8'hFF;
            14'd4751: data <= 8'hFF;
            14'd4752: data <= 8'hFF;
            14'd4753: data <= 8'hF0;
            14'd4754: data <= 8'h00;
            14'd4755: data <= 8'h00;
            14'd4756: data <= 8'h00;
            14'd4757: data <= 8'h00;
            14'd4758: data <= 8'h00;
            14'd4759: data <= 8'h00;
            14'd4760: data <= 8'h00;
            14'd4761: data <= 8'h00;
            14'd4762: data <= 8'h00;
            14'd4763: data <= 8'h00;
            14'd4764: data <= 8'h00;
            14'd4765: data <= 8'h00;
            14'd4766: data <= 8'h0F;
            14'd4767: data <= 8'hFF;
            14'd4768: data <= 8'hFF;
            14'd4769: data <= 8'hFF;
            14'd4770: data <= 8'hFF;
            14'd4771: data <= 8'hFF;
            14'd4772: data <= 8'hFF;
            14'd4773: data <= 8'hFF;
            14'd4774: data <= 8'hFF;
            14'd4775: data <= 8'hFF;
            14'd4776: data <= 8'hFF;
            14'd4777: data <= 8'hFF;
            14'd4778: data <= 8'hFF;
            14'd4779: data <= 8'hFF;
            14'd4780: data <= 8'hFF;
            14'd4781: data <= 8'hFF;
            14'd4782: data <= 8'hE0;
            14'd4783: data <= 8'h3F;
            14'd4784: data <= 8'hFC;
            14'd4785: data <= 8'h07;
            14'd4786: data <= 8'hFF;
            14'd4787: data <= 8'hFF;
            14'd4788: data <= 8'hFF;
            14'd4789: data <= 8'hFF;
            14'd4790: data <= 8'hFF;
            14'd4791: data <= 8'hFF;
            14'd4792: data <= 8'hFF;
            14'd4793: data <= 8'hF0;
            14'd4794: data <= 8'h00;
            14'd4795: data <= 8'h00;
            14'd4796: data <= 8'h00;
            14'd4797: data <= 8'h00;
            14'd4798: data <= 8'h00;
            14'd4799: data <= 8'h00;
            14'd4800: data <= 8'h00;
            14'd4801: data <= 8'h00;
            14'd4802: data <= 8'h00;
            14'd4803: data <= 8'h00;
            14'd4804: data <= 8'h00;
            14'd4805: data <= 8'h00;
            14'd4806: data <= 8'h0F;
            14'd4807: data <= 8'hFF;
            14'd4808: data <= 8'hFF;
            14'd4809: data <= 8'hFF;
            14'd4810: data <= 8'hFF;
            14'd4811: data <= 8'hFF;
            14'd4812: data <= 8'hFF;
            14'd4813: data <= 8'hFF;
            14'd4814: data <= 8'hFF;
            14'd4815: data <= 8'hFF;
            14'd4816: data <= 8'hFF;
            14'd4817: data <= 8'hFF;
            14'd4818: data <= 8'hFF;
            14'd4819: data <= 8'hFF;
            14'd4820: data <= 8'hFF;
            14'd4821: data <= 8'hFF;
            14'd4822: data <= 8'hE0;
            14'd4823: data <= 8'h77;
            14'd4824: data <= 8'hF8;
            14'd4825: data <= 8'h0F;
            14'd4826: data <= 8'hFF;
            14'd4827: data <= 8'hFF;
            14'd4828: data <= 8'hFF;
            14'd4829: data <= 8'hFF;
            14'd4830: data <= 8'hFF;
            14'd4831: data <= 8'hFF;
            14'd4832: data <= 8'hFF;
            14'd4833: data <= 8'hF0;
            14'd4834: data <= 8'h00;
            14'd4835: data <= 8'h00;
            14'd4836: data <= 8'h00;
            14'd4837: data <= 8'h00;
            14'd4838: data <= 8'h00;
            14'd4839: data <= 8'h00;
            14'd4840: data <= 8'h00;
            14'd4841: data <= 8'h00;
            14'd4842: data <= 8'h00;
            14'd4843: data <= 8'h00;
            14'd4844: data <= 8'h00;
            14'd4845: data <= 8'h00;
            14'd4846: data <= 8'h0F;
            14'd4847: data <= 8'hFF;
            14'd4848: data <= 8'hFF;
            14'd4849: data <= 8'hFF;
            14'd4850: data <= 8'hFF;
            14'd4851: data <= 8'hFF;
            14'd4852: data <= 8'hFF;
            14'd4853: data <= 8'hFF;
            14'd4854: data <= 8'hFF;
            14'd4855: data <= 8'hFF;
            14'd4856: data <= 8'hFF;
            14'd4857: data <= 8'hFF;
            14'd4858: data <= 8'hFF;
            14'd4859: data <= 8'hFF;
            14'd4860: data <= 8'hFF;
            14'd4861: data <= 8'hFF;
            14'd4862: data <= 8'hE0;
            14'd4863: data <= 8'h7F;
            14'd4864: data <= 8'hF0;
            14'd4865: data <= 8'h1F;
            14'd4866: data <= 8'hFF;
            14'd4867: data <= 8'hFF;
            14'd4868: data <= 8'hFF;
            14'd4869: data <= 8'hFF;
            14'd4870: data <= 8'hFF;
            14'd4871: data <= 8'hFF;
            14'd4872: data <= 8'hFF;
            14'd4873: data <= 8'hF0;
            14'd4874: data <= 8'h00;
            14'd4875: data <= 8'h00;
            14'd4876: data <= 8'h00;
            14'd4877: data <= 8'h00;
            14'd4878: data <= 8'h00;
            14'd4879: data <= 8'h00;
            14'd4880: data <= 8'h00;
            14'd4881: data <= 8'h00;
            14'd4882: data <= 8'h00;
            14'd4883: data <= 8'h00;
            14'd4884: data <= 8'h00;
            14'd4885: data <= 8'h00;
            14'd4886: data <= 8'h0F;
            14'd4887: data <= 8'hFF;
            14'd4888: data <= 8'hFF;
            14'd4889: data <= 8'hFF;
            14'd4890: data <= 8'hFF;
            14'd4891: data <= 8'hFF;
            14'd4892: data <= 8'hFF;
            14'd4893: data <= 8'hFF;
            14'd4894: data <= 8'hDF;
            14'd4895: data <= 8'hFF;
            14'd4896: data <= 8'hFF;
            14'd4897: data <= 8'hFF;
            14'd4898: data <= 8'hFF;
            14'd4899: data <= 8'hFF;
            14'd4900: data <= 8'hFF;
            14'd4901: data <= 8'hFF;
            14'd4902: data <= 8'hE0;
            14'd4903: data <= 8'hFF;
            14'd4904: data <= 8'hE0;
            14'd4905: data <= 8'h1F;
            14'd4906: data <= 8'hFF;
            14'd4907: data <= 8'hFF;
            14'd4908: data <= 8'hFF;
            14'd4909: data <= 8'hFF;
            14'd4910: data <= 8'hFF;
            14'd4911: data <= 8'hBF;
            14'd4912: data <= 8'hFF;
            14'd4913: data <= 8'hF0;
            14'd4914: data <= 8'h00;
            14'd4915: data <= 8'h00;
            14'd4916: data <= 8'h00;
            14'd4917: data <= 8'h00;
            14'd4918: data <= 8'h00;
            14'd4919: data <= 8'h00;
            14'd4920: data <= 8'h00;
            14'd4921: data <= 8'h00;
            14'd4922: data <= 8'h00;
            14'd4923: data <= 8'h00;
            14'd4924: data <= 8'h00;
            14'd4925: data <= 8'h00;
            14'd4926: data <= 8'h0F;
            14'd4927: data <= 8'hFF;
            14'd4928: data <= 8'hFF;
            14'd4929: data <= 8'hFF;
            14'd4930: data <= 8'hFF;
            14'd4931: data <= 8'hFF;
            14'd4932: data <= 8'hFF;
            14'd4933: data <= 8'hFF;
            14'd4934: data <= 8'hFF;
            14'd4935: data <= 8'hFF;
            14'd4936: data <= 8'hFF;
            14'd4937: data <= 8'hFF;
            14'd4938: data <= 8'hFF;
            14'd4939: data <= 8'hFF;
            14'd4940: data <= 8'hFF;
            14'd4941: data <= 8'hFF;
            14'd4942: data <= 8'hC0;
            14'd4943: data <= 8'hFF;
            14'd4944: data <= 8'hC0;
            14'd4945: data <= 8'h3F;
            14'd4946: data <= 8'hFF;
            14'd4947: data <= 8'hFF;
            14'd4948: data <= 8'hFF;
            14'd4949: data <= 8'hFF;
            14'd4950: data <= 8'hFF;
            14'd4951: data <= 8'hFF;
            14'd4952: data <= 8'hFF;
            14'd4953: data <= 8'hF0;
            14'd4954: data <= 8'h00;
            14'd4955: data <= 8'h00;
            14'd4956: data <= 8'h00;
            14'd4957: data <= 8'h00;
            14'd4958: data <= 8'h00;
            14'd4959: data <= 8'h00;
            14'd4960: data <= 8'h00;
            14'd4961: data <= 8'h00;
            14'd4962: data <= 8'h00;
            14'd4963: data <= 8'h00;
            14'd4964: data <= 8'h00;
            14'd4965: data <= 8'h00;
            14'd4966: data <= 8'h0F;
            14'd4967: data <= 8'hFF;
            14'd4968: data <= 8'hFF;
            14'd4969: data <= 8'hFF;
            14'd4970: data <= 8'hFF;
            14'd4971: data <= 8'hFF;
            14'd4972: data <= 8'hFF;
            14'd4973: data <= 8'hFF;
            14'd4974: data <= 8'hFF;
            14'd4975: data <= 8'hFF;
            14'd4976: data <= 8'hFF;
            14'd4977: data <= 8'hFF;
            14'd4978: data <= 8'hFF;
            14'd4979: data <= 8'hFF;
            14'd4980: data <= 8'hFF;
            14'd4981: data <= 8'hFF;
            14'd4982: data <= 8'hC1;
            14'd4983: data <= 8'hFF;
            14'd4984: data <= 8'h80;
            14'd4985: data <= 8'h7F;
            14'd4986: data <= 8'hFF;
            14'd4987: data <= 8'hFF;
            14'd4988: data <= 8'hFF;
            14'd4989: data <= 8'hFF;
            14'd4990: data <= 8'hFF;
            14'd4991: data <= 8'hFF;
            14'd4992: data <= 8'hFF;
            14'd4993: data <= 8'hF0;
            14'd4994: data <= 8'h00;
            14'd4995: data <= 8'h00;
            14'd4996: data <= 8'h00;
            14'd4997: data <= 8'h00;
            14'd4998: data <= 8'h00;
            14'd4999: data <= 8'h00;
            14'd5000: data <= 8'h00;
            14'd5001: data <= 8'h00;
            14'd5002: data <= 8'h00;
            14'd5003: data <= 8'h00;
            14'd5004: data <= 8'h00;
            14'd5005: data <= 8'h00;
            14'd5006: data <= 8'h0F;
            14'd5007: data <= 8'hFF;
            14'd5008: data <= 8'hFF;
            14'd5009: data <= 8'hFF;
            14'd5010: data <= 8'hFF;
            14'd5011: data <= 8'hFF;
            14'd5012: data <= 8'hFF;
            14'd5013: data <= 8'hFF;
            14'd5014: data <= 8'hFF;
            14'd5015: data <= 8'hFF;
            14'd5016: data <= 8'hFF;
            14'd5017: data <= 8'hFF;
            14'd5018: data <= 8'hFF;
            14'd5019: data <= 8'hFF;
            14'd5020: data <= 8'hFF;
            14'd5021: data <= 8'hFF;
            14'd5022: data <= 8'hC1;
            14'd5023: data <= 8'hFF;
            14'd5024: data <= 8'h00;
            14'd5025: data <= 8'h7F;
            14'd5026: data <= 8'hFF;
            14'd5027: data <= 8'hFF;
            14'd5028: data <= 8'hFF;
            14'd5029: data <= 8'hFF;
            14'd5030: data <= 8'hFF;
            14'd5031: data <= 8'hFF;
            14'd5032: data <= 8'hFF;
            14'd5033: data <= 8'hF0;
            14'd5034: data <= 8'h00;
            14'd5035: data <= 8'h00;
            14'd5036: data <= 8'h00;
            14'd5037: data <= 8'h00;
            14'd5038: data <= 8'h00;
            14'd5039: data <= 8'h00;
            14'd5040: data <= 8'h00;
            14'd5041: data <= 8'h00;
            14'd5042: data <= 8'h00;
            14'd5043: data <= 8'h00;
            14'd5044: data <= 8'h00;
            14'd5045: data <= 8'h00;
            14'd5046: data <= 8'h0F;
            14'd5047: data <= 8'hFF;
            14'd5048: data <= 8'hFF;
            14'd5049: data <= 8'hFF;
            14'd5050: data <= 8'hFF;
            14'd5051: data <= 8'hFF;
            14'd5052: data <= 8'hFF;
            14'd5053: data <= 8'hFF;
            14'd5054: data <= 8'hFF;
            14'd5055: data <= 8'hFF;
            14'd5056: data <= 8'hFF;
            14'd5057: data <= 8'hFF;
            14'd5058: data <= 8'hFF;
            14'd5059: data <= 8'hFF;
            14'd5060: data <= 8'hFF;
            14'd5061: data <= 8'hFF;
            14'd5062: data <= 8'hC1;
            14'd5063: data <= 8'hFE;
            14'd5064: data <= 8'h01;
            14'd5065: data <= 8'hFF;
            14'd5066: data <= 8'hFF;
            14'd5067: data <= 8'hFF;
            14'd5068: data <= 8'hFF;
            14'd5069: data <= 8'hFF;
            14'd5070: data <= 8'hFF;
            14'd5071: data <= 8'hFF;
            14'd5072: data <= 8'hFF;
            14'd5073: data <= 8'hF0;
            14'd5074: data <= 8'h00;
            14'd5075: data <= 8'h00;
            14'd5076: data <= 8'h00;
            14'd5077: data <= 8'h00;
            14'd5078: data <= 8'h00;
            14'd5079: data <= 8'h00;
            14'd5080: data <= 8'h00;
            14'd5081: data <= 8'h00;
            14'd5082: data <= 8'h00;
            14'd5083: data <= 8'h00;
            14'd5084: data <= 8'h00;
            14'd5085: data <= 8'h00;
            14'd5086: data <= 8'h0F;
            14'd5087: data <= 8'hFF;
            14'd5088: data <= 8'hFF;
            14'd5089: data <= 8'hFF;
            14'd5090: data <= 8'hFF;
            14'd5091: data <= 8'hFF;
            14'd5092: data <= 8'hFF;
            14'd5093: data <= 8'hFF;
            14'd5094: data <= 8'hFF;
            14'd5095: data <= 8'hFF;
            14'd5096: data <= 8'hFF;
            14'd5097: data <= 8'hFF;
            14'd5098: data <= 8'hFF;
            14'd5099: data <= 8'hFF;
            14'd5100: data <= 8'hFF;
            14'd5101: data <= 8'hFF;
            14'd5102: data <= 8'h83;
            14'd5103: data <= 8'hFC;
            14'd5104: data <= 8'h01;
            14'd5105: data <= 8'hFF;
            14'd5106: data <= 8'hFF;
            14'd5107: data <= 8'hFF;
            14'd5108: data <= 8'hFF;
            14'd5109: data <= 8'hFF;
            14'd5110: data <= 8'hFF;
            14'd5111: data <= 8'hFF;
            14'd5112: data <= 8'hFF;
            14'd5113: data <= 8'hF0;
            14'd5114: data <= 8'h00;
            14'd5115: data <= 8'h00;
            14'd5116: data <= 8'h00;
            14'd5117: data <= 8'h00;
            14'd5118: data <= 8'h00;
            14'd5119: data <= 8'h00;
            14'd5120: data <= 8'h00;
            14'd5121: data <= 8'h00;
            14'd5122: data <= 8'h00;
            14'd5123: data <= 8'h00;
            14'd5124: data <= 8'h00;
            14'd5125: data <= 8'h00;
            14'd5126: data <= 8'h0F;
            14'd5127: data <= 8'hFF;
            14'd5128: data <= 8'hFF;
            14'd5129: data <= 8'hFF;
            14'd5130: data <= 8'hFE;
            14'd5131: data <= 8'hFF;
            14'd5132: data <= 8'hFF;
            14'd5133: data <= 8'hFF;
            14'd5134: data <= 8'hFF;
            14'd5135: data <= 8'hFF;
            14'd5136: data <= 8'hFF;
            14'd5137: data <= 8'hFF;
            14'd5138: data <= 8'hFF;
            14'd5139: data <= 8'hFF;
            14'd5140: data <= 8'hFF;
            14'd5141: data <= 8'hFF;
            14'd5142: data <= 8'hC3;
            14'd5143: data <= 8'hF8;
            14'd5144: data <= 8'h07;
            14'd5145: data <= 8'hFF;
            14'd5146: data <= 8'hFF;
            14'd5147: data <= 8'hFF;
            14'd5148: data <= 8'hFF;
            14'd5149: data <= 8'hFF;
            14'd5150: data <= 8'hFF;
            14'd5151: data <= 8'hFF;
            14'd5152: data <= 8'hFF;
            14'd5153: data <= 8'hF0;
            14'd5154: data <= 8'h00;
            14'd5155: data <= 8'h00;
            14'd5156: data <= 8'h00;
            14'd5157: data <= 8'h00;
            14'd5158: data <= 8'h00;
            14'd5159: data <= 8'h00;
            14'd5160: data <= 8'h00;
            14'd5161: data <= 8'h00;
            14'd5162: data <= 8'h00;
            14'd5163: data <= 8'h00;
            14'd5164: data <= 8'h00;
            14'd5165: data <= 8'h00;
            14'd5166: data <= 8'h0F;
            14'd5167: data <= 8'hFF;
            14'd5168: data <= 8'hFF;
            14'd5169: data <= 8'hFF;
            14'd5170: data <= 8'hFF;
            14'd5171: data <= 8'hBF;
            14'd5172: data <= 8'hFF;
            14'd5173: data <= 8'hFF;
            14'd5174: data <= 8'hFF;
            14'd5175: data <= 8'hFF;
            14'd5176: data <= 8'hFF;
            14'd5177: data <= 8'hFF;
            14'd5178: data <= 8'hFF;
            14'd5179: data <= 8'hFF;
            14'd5180: data <= 8'hFF;
            14'd5181: data <= 8'hFF;
            14'd5182: data <= 8'h83;
            14'd5183: data <= 8'hF0;
            14'd5184: data <= 8'h06;
            14'd5185: data <= 8'hFF;
            14'd5186: data <= 8'hFF;
            14'd5187: data <= 8'hFF;
            14'd5188: data <= 8'hFF;
            14'd5189: data <= 8'hFB;
            14'd5190: data <= 8'hFF;
            14'd5191: data <= 8'hFF;
            14'd5192: data <= 8'hFF;
            14'd5193: data <= 8'hF0;
            14'd5194: data <= 8'h00;
            14'd5195: data <= 8'h00;
            14'd5196: data <= 8'h00;
            14'd5197: data <= 8'h00;
            14'd5198: data <= 8'h00;
            14'd5199: data <= 8'h00;
            14'd5200: data <= 8'h00;
            14'd5201: data <= 8'h00;
            14'd5202: data <= 8'h00;
            14'd5203: data <= 8'h00;
            14'd5204: data <= 8'h00;
            14'd5205: data <= 8'h00;
            14'd5206: data <= 8'h0F;
            14'd5207: data <= 8'hFF;
            14'd5208: data <= 8'hFF;
            14'd5209: data <= 8'hFF;
            14'd5210: data <= 8'hFF;
            14'd5211: data <= 8'hFF;
            14'd5212: data <= 8'hFF;
            14'd5213: data <= 8'hFF;
            14'd5214: data <= 8'hFF;
            14'd5215: data <= 8'hFF;
            14'd5216: data <= 8'hFF;
            14'd5217: data <= 8'hFF;
            14'd5218: data <= 8'hFF;
            14'd5219: data <= 8'hFF;
            14'd5220: data <= 8'hFF;
            14'd5221: data <= 8'hFF;
            14'd5222: data <= 8'h83;
            14'd5223: data <= 8'hC0;
            14'd5224: data <= 8'h0F;
            14'd5225: data <= 8'hFF;
            14'd5226: data <= 8'hFF;
            14'd5227: data <= 8'hFF;
            14'd5228: data <= 8'hFF;
            14'd5229: data <= 8'hFF;
            14'd5230: data <= 8'hFF;
            14'd5231: data <= 8'hFF;
            14'd5232: data <= 8'hFF;
            14'd5233: data <= 8'hF0;
            14'd5234: data <= 8'h00;
            14'd5235: data <= 8'h00;
            14'd5236: data <= 8'h00;
            14'd5237: data <= 8'h00;
            14'd5238: data <= 8'h00;
            14'd5239: data <= 8'h00;
            14'd5240: data <= 8'h00;
            14'd5241: data <= 8'h00;
            14'd5242: data <= 8'h00;
            14'd5243: data <= 8'h00;
            14'd5244: data <= 8'h00;
            14'd5245: data <= 8'h00;
            14'd5246: data <= 8'h0F;
            14'd5247: data <= 8'hFF;
            14'd5248: data <= 8'hFF;
            14'd5249: data <= 8'hFF;
            14'd5250: data <= 8'hFF;
            14'd5251: data <= 8'hFF;
            14'd5252: data <= 8'hFF;
            14'd5253: data <= 8'hFF;
            14'd5254: data <= 8'hFF;
            14'd5255: data <= 8'hFF;
            14'd5256: data <= 8'hFF;
            14'd5257: data <= 8'hFF;
            14'd5258: data <= 8'hFF;
            14'd5259: data <= 8'hFF;
            14'd5260: data <= 8'hFF;
            14'd5261: data <= 8'hFF;
            14'd5262: data <= 8'h81;
            14'd5263: data <= 8'h00;
            14'd5264: data <= 8'h1F;
            14'd5265: data <= 8'hFF;
            14'd5266: data <= 8'hFF;
            14'd5267: data <= 8'hFF;
            14'd5268: data <= 8'hFF;
            14'd5269: data <= 8'hFF;
            14'd5270: data <= 8'hFF;
            14'd5271: data <= 8'hFF;
            14'd5272: data <= 8'hFF;
            14'd5273: data <= 8'hF0;
            14'd5274: data <= 8'h00;
            14'd5275: data <= 8'h00;
            14'd5276: data <= 8'h00;
            14'd5277: data <= 8'h00;
            14'd5278: data <= 8'h00;
            14'd5279: data <= 8'h00;
            14'd5280: data <= 8'h00;
            14'd5281: data <= 8'h00;
            14'd5282: data <= 8'h00;
            14'd5283: data <= 8'h00;
            14'd5284: data <= 8'h00;
            14'd5285: data <= 8'h00;
            14'd5286: data <= 8'h0F;
            14'd5287: data <= 8'hFF;
            14'd5288: data <= 8'hFF;
            14'd5289: data <= 8'hFF;
            14'd5290: data <= 8'hFF;
            14'd5291: data <= 8'hFF;
            14'd5292: data <= 8'hFF;
            14'd5293: data <= 8'hFF;
            14'd5294: data <= 8'hFF;
            14'd5295: data <= 8'hFF;
            14'd5296: data <= 8'hFF;
            14'd5297: data <= 8'hFF;
            14'd5298: data <= 8'hFF;
            14'd5299: data <= 8'hFF;
            14'd5300: data <= 8'hFF;
            14'd5301: data <= 8'hFF;
            14'd5302: data <= 8'h80;
            14'd5303: data <= 8'h00;
            14'd5304: data <= 8'h3F;
            14'd5305: data <= 8'hFF;
            14'd5306: data <= 8'hFF;
            14'd5307: data <= 8'hFF;
            14'd5308: data <= 8'hFF;
            14'd5309: data <= 8'hFF;
            14'd5310: data <= 8'hFF;
            14'd5311: data <= 8'hFF;
            14'd5312: data <= 8'hFF;
            14'd5313: data <= 8'hF0;
            14'd5314: data <= 8'h00;
            14'd5315: data <= 8'h00;
            14'd5316: data <= 8'h00;
            14'd5317: data <= 8'h00;
            14'd5318: data <= 8'h00;
            14'd5319: data <= 8'h00;
            14'd5320: data <= 8'h00;
            14'd5321: data <= 8'h00;
            14'd5322: data <= 8'h00;
            14'd5323: data <= 8'h00;
            14'd5324: data <= 8'h00;
            14'd5325: data <= 8'h00;
            14'd5326: data <= 8'h0F;
            14'd5327: data <= 8'hFF;
            14'd5328: data <= 8'hFF;
            14'd5329: data <= 8'hFF;
            14'd5330: data <= 8'hFF;
            14'd5331: data <= 8'hFF;
            14'd5332: data <= 8'hFF;
            14'd5333: data <= 8'hFF;
            14'd5334: data <= 8'hFF;
            14'd5335: data <= 8'hFF;
            14'd5336: data <= 8'hFF;
            14'd5337: data <= 8'hFF;
            14'd5338: data <= 8'hFF;
            14'd5339: data <= 8'hFF;
            14'd5340: data <= 8'hFF;
            14'd5341: data <= 8'hFF;
            14'd5342: data <= 8'hC0;
            14'd5343: data <= 8'h00;
            14'd5344: data <= 8'h7F;
            14'd5345: data <= 8'hFF;
            14'd5346: data <= 8'hFF;
            14'd5347: data <= 8'hFF;
            14'd5348: data <= 8'hFF;
            14'd5349: data <= 8'hFF;
            14'd5350: data <= 8'hFF;
            14'd5351: data <= 8'hFF;
            14'd5352: data <= 8'hFF;
            14'd5353: data <= 8'hF0;
            14'd5354: data <= 8'h00;
            14'd5355: data <= 8'h00;
            14'd5356: data <= 8'h00;
            14'd5357: data <= 8'h00;
            14'd5358: data <= 8'h00;
            14'd5359: data <= 8'h00;
            14'd5360: data <= 8'h00;
            14'd5361: data <= 8'h00;
            14'd5362: data <= 8'h00;
            14'd5363: data <= 8'h00;
            14'd5364: data <= 8'h00;
            14'd5365: data <= 8'h00;
            14'd5366: data <= 8'h0F;
            14'd5367: data <= 8'hFF;
            14'd5368: data <= 8'hFF;
            14'd5369: data <= 8'hFF;
            14'd5370: data <= 8'hFF;
            14'd5371: data <= 8'hFF;
            14'd5372: data <= 8'hFF;
            14'd5373: data <= 8'hFF;
            14'd5374: data <= 8'hFF;
            14'd5375: data <= 8'hFF;
            14'd5376: data <= 8'hFF;
            14'd5377: data <= 8'hFF;
            14'd5378: data <= 8'hFF;
            14'd5379: data <= 8'hFF;
            14'd5380: data <= 8'hFF;
            14'd5381: data <= 8'hFF;
            14'd5382: data <= 8'h40;
            14'd5383: data <= 8'h01;
            14'd5384: data <= 8'hFF;
            14'd5385: data <= 8'hFF;
            14'd5386: data <= 8'hFF;
            14'd5387: data <= 8'hFF;
            14'd5388: data <= 8'hFF;
            14'd5389: data <= 8'hFF;
            14'd5390: data <= 8'hFF;
            14'd5391: data <= 8'hFF;
            14'd5392: data <= 8'hFF;
            14'd5393: data <= 8'hF0;
            14'd5394: data <= 8'h00;
            14'd5395: data <= 8'h00;
            14'd5396: data <= 8'h00;
            14'd5397: data <= 8'h00;
            14'd5398: data <= 8'h00;
            14'd5399: data <= 8'h00;
            14'd5400: data <= 8'h00;
            14'd5401: data <= 8'h00;
            14'd5402: data <= 8'h00;
            14'd5403: data <= 8'h00;
            14'd5404: data <= 8'h00;
            14'd5405: data <= 8'h00;
            14'd5406: data <= 8'h0F;
            14'd5407: data <= 8'hFF;
            14'd5408: data <= 8'hFF;
            14'd5409: data <= 8'hFF;
            14'd5410: data <= 8'hFF;
            14'd5411: data <= 8'hFF;
            14'd5412: data <= 8'hFF;
            14'd5413: data <= 8'hFF;
            14'd5414: data <= 8'hFF;
            14'd5415: data <= 8'hFF;
            14'd5416: data <= 8'hFF;
            14'd5417: data <= 8'hFF;
            14'd5418: data <= 8'hFF;
            14'd5419: data <= 8'hFF;
            14'd5420: data <= 8'hE7;
            14'd5421: data <= 8'hFF;
            14'd5422: data <= 8'hE0;
            14'd5423: data <= 8'h07;
            14'd5424: data <= 8'hFF;
            14'd5425: data <= 8'hFF;
            14'd5426: data <= 8'hFF;
            14'd5427: data <= 8'hFF;
            14'd5428: data <= 8'hFF;
            14'd5429: data <= 8'hFF;
            14'd5430: data <= 8'hFF;
            14'd5431: data <= 8'hFF;
            14'd5432: data <= 8'hFF;
            14'd5433: data <= 8'hF0;
            14'd5434: data <= 8'h00;
            14'd5435: data <= 8'h00;
            14'd5436: data <= 8'h00;
            14'd5437: data <= 8'h00;
            14'd5438: data <= 8'h00;
            14'd5439: data <= 8'h00;
            14'd5440: data <= 8'h00;
            14'd5441: data <= 8'h00;
            14'd5442: data <= 8'h00;
            14'd5443: data <= 8'h00;
            14'd5444: data <= 8'h00;
            14'd5445: data <= 8'h00;
            14'd5446: data <= 8'h0F;
            14'd5447: data <= 8'hFF;
            14'd5448: data <= 8'hFF;
            14'd5449: data <= 8'hFF;
            14'd5450: data <= 8'hFF;
            14'd5451: data <= 8'hFF;
            14'd5452: data <= 8'hFF;
            14'd5453: data <= 8'hFF;
            14'd5454: data <= 8'hFF;
            14'd5455: data <= 8'hFF;
            14'd5456: data <= 8'hFF;
            14'd5457: data <= 8'hFF;
            14'd5458: data <= 8'hFF;
            14'd5459: data <= 8'hFF;
            14'd5460: data <= 8'hC3;
            14'd5461: data <= 8'h7F;
            14'd5462: data <= 8'hF0;
            14'd5463: data <= 8'h1F;
            14'd5464: data <= 8'hFF;
            14'd5465: data <= 8'hFF;
            14'd5466: data <= 8'hFF;
            14'd5467: data <= 8'hFF;
            14'd5468: data <= 8'hFF;
            14'd5469: data <= 8'hFF;
            14'd5470: data <= 8'hFF;
            14'd5471: data <= 8'hFF;
            14'd5472: data <= 8'hFF;
            14'd5473: data <= 8'hF0;
            14'd5474: data <= 8'h00;
            14'd5475: data <= 8'h00;
            14'd5476: data <= 8'h00;
            14'd5477: data <= 8'h00;
            14'd5478: data <= 8'h00;
            14'd5479: data <= 8'h00;
            14'd5480: data <= 8'h00;
            14'd5481: data <= 8'h00;
            14'd5482: data <= 8'h00;
            14'd5483: data <= 8'h00;
            14'd5484: data <= 8'h00;
            14'd5485: data <= 8'h00;
            14'd5486: data <= 8'h0F;
            14'd5487: data <= 8'hFF;
            14'd5488: data <= 8'hFF;
            14'd5489: data <= 8'hFF;
            14'd5490: data <= 8'hFF;
            14'd5491: data <= 8'hFF;
            14'd5492: data <= 8'hFF;
            14'd5493: data <= 8'hFF;
            14'd5494: data <= 8'hFF;
            14'd5495: data <= 8'hFF;
            14'd5496: data <= 8'hFF;
            14'd5497: data <= 8'hFF;
            14'd5498: data <= 8'hFF;
            14'd5499: data <= 8'hFF;
            14'd5500: data <= 8'h87;
            14'd5501: data <= 8'hFF;
            14'd5502: data <= 8'hFF;
            14'd5503: data <= 8'hFB;
            14'd5504: data <= 8'hFF;
            14'd5505: data <= 8'hFF;
            14'd5506: data <= 8'hFF;
            14'd5507: data <= 8'hFF;
            14'd5508: data <= 8'hFF;
            14'd5509: data <= 8'hFF;
            14'd5510: data <= 8'hFF;
            14'd5511: data <= 8'hFF;
            14'd5512: data <= 8'hFF;
            14'd5513: data <= 8'hF0;
            14'd5514: data <= 8'h00;
            14'd5515: data <= 8'h00;
            14'd5516: data <= 8'h00;
            14'd5517: data <= 8'h00;
            14'd5518: data <= 8'h00;
            14'd5519: data <= 8'h00;
            14'd5520: data <= 8'h00;
            14'd5521: data <= 8'h00;
            14'd5522: data <= 8'h00;
            14'd5523: data <= 8'h00;
            14'd5524: data <= 8'h00;
            14'd5525: data <= 8'h00;
            14'd5526: data <= 8'h0F;
            14'd5527: data <= 8'hFF;
            14'd5528: data <= 8'hFF;
            14'd5529: data <= 8'hFF;
            14'd5530: data <= 8'hFF;
            14'd5531: data <= 8'hFF;
            14'd5532: data <= 8'hFF;
            14'd5533: data <= 8'hFF;
            14'd5534: data <= 8'hFF;
            14'd5535: data <= 8'hFF;
            14'd5536: data <= 8'hFF;
            14'd5537: data <= 8'hFF;
            14'd5538: data <= 8'hFF;
            14'd5539: data <= 8'hFF;
            14'd5540: data <= 8'h07;
            14'd5541: data <= 8'hFF;
            14'd5542: data <= 8'hFF;
            14'd5543: data <= 8'hFF;
            14'd5544: data <= 8'hFF;
            14'd5545: data <= 8'hFF;
            14'd5546: data <= 8'hFF;
            14'd5547: data <= 8'hFF;
            14'd5548: data <= 8'hFF;
            14'd5549: data <= 8'hFF;
            14'd5550: data <= 8'hFF;
            14'd5551: data <= 8'hFF;
            14'd5552: data <= 8'hFF;
            14'd5553: data <= 8'hF0;
            14'd5554: data <= 8'h00;
            14'd5555: data <= 8'h00;
            14'd5556: data <= 8'h00;
            14'd5557: data <= 8'h00;
            14'd5558: data <= 8'h00;
            14'd5559: data <= 8'h00;
            14'd5560: data <= 8'h00;
            14'd5561: data <= 8'h00;
            14'd5562: data <= 8'h00;
            14'd5563: data <= 8'h00;
            14'd5564: data <= 8'h00;
            14'd5565: data <= 8'h00;
            14'd5566: data <= 8'h0F;
            14'd5567: data <= 8'hFF;
            14'd5568: data <= 8'hFF;
            14'd5569: data <= 8'hFF;
            14'd5570: data <= 8'hFF;
            14'd5571: data <= 8'hFF;
            14'd5572: data <= 8'hFF;
            14'd5573: data <= 8'hFF;
            14'd5574: data <= 8'hFF;
            14'd5575: data <= 8'hFF;
            14'd5576: data <= 8'hFF;
            14'd5577: data <= 8'hFF;
            14'd5578: data <= 8'hFF;
            14'd5579: data <= 8'hFF;
            14'd5580: data <= 8'h0F;
            14'd5581: data <= 8'hCF;
            14'd5582: data <= 8'hFF;
            14'd5583: data <= 8'hFF;
            14'd5584: data <= 8'hFF;
            14'd5585: data <= 8'hFF;
            14'd5586: data <= 8'hFF;
            14'd5587: data <= 8'hFF;
            14'd5588: data <= 8'hFF;
            14'd5589: data <= 8'hFF;
            14'd5590: data <= 8'hFF;
            14'd5591: data <= 8'hFF;
            14'd5592: data <= 8'hFF;
            14'd5593: data <= 8'hF0;
            14'd5594: data <= 8'h00;
            14'd5595: data <= 8'h00;
            14'd5596: data <= 8'h00;
            14'd5597: data <= 8'h00;
            14'd5598: data <= 8'h00;
            14'd5599: data <= 8'h00;
            14'd5600: data <= 8'h00;
            14'd5601: data <= 8'h00;
            14'd5602: data <= 8'h00;
            14'd5603: data <= 8'h00;
            14'd5604: data <= 8'h00;
            14'd5605: data <= 8'h00;
            14'd5606: data <= 8'h0F;
            14'd5607: data <= 8'hFF;
            14'd5608: data <= 8'hFF;
            14'd5609: data <= 8'hFF;
            14'd5610: data <= 8'hFF;
            14'd5611: data <= 8'hFF;
            14'd5612: data <= 8'hFF;
            14'd5613: data <= 8'hFF;
            14'd5614: data <= 8'hFF;
            14'd5615: data <= 8'hFF;
            14'd5616: data <= 8'hFF;
            14'd5617: data <= 8'hFF;
            14'd5618: data <= 8'hFF;
            14'd5619: data <= 8'hFE;
            14'd5620: data <= 8'h1F;
            14'd5621: data <= 8'h87;
            14'd5622: data <= 8'hFE;
            14'd5623: data <= 8'h7F;
            14'd5624: data <= 8'hFF;
            14'd5625: data <= 8'hFF;
            14'd5626: data <= 8'hFF;
            14'd5627: data <= 8'hFF;
            14'd5628: data <= 8'hFF;
            14'd5629: data <= 8'hFF;
            14'd5630: data <= 8'hFF;
            14'd5631: data <= 8'hFF;
            14'd5632: data <= 8'hFF;
            14'd5633: data <= 8'hF0;
            14'd5634: data <= 8'h00;
            14'd5635: data <= 8'h00;
            14'd5636: data <= 8'h00;
            14'd5637: data <= 8'h00;
            14'd5638: data <= 8'h00;
            14'd5639: data <= 8'h00;
            14'd5640: data <= 8'h00;
            14'd5641: data <= 8'h00;
            14'd5642: data <= 8'h00;
            14'd5643: data <= 8'h00;
            14'd5644: data <= 8'h00;
            14'd5645: data <= 8'h00;
            14'd5646: data <= 8'h0F;
            14'd5647: data <= 8'hFF;
            14'd5648: data <= 8'hFF;
            14'd5649: data <= 8'hFF;
            14'd5650: data <= 8'hFF;
            14'd5651: data <= 8'hFF;
            14'd5652: data <= 8'hFF;
            14'd5653: data <= 8'hFF;
            14'd5654: data <= 8'hFF;
            14'd5655: data <= 8'hFF;
            14'd5656: data <= 8'hFF;
            14'd5657: data <= 8'hFF;
            14'd5658: data <= 8'hFF;
            14'd5659: data <= 8'hFC;
            14'd5660: data <= 8'h1F;
            14'd5661: data <= 8'h87;
            14'd5662: data <= 8'hFC;
            14'd5663: data <= 8'h3F;
            14'd5664: data <= 8'hFF;
            14'd5665: data <= 8'hFF;
            14'd5666: data <= 8'hFF;
            14'd5667: data <= 8'hFF;
            14'd5668: data <= 8'hFF;
            14'd5669: data <= 8'hFF;
            14'd5670: data <= 8'hFF;
            14'd5671: data <= 8'hFF;
            14'd5672: data <= 8'hFF;
            14'd5673: data <= 8'hF0;
            14'd5674: data <= 8'h00;
            14'd5675: data <= 8'h00;
            14'd5676: data <= 8'h00;
            14'd5677: data <= 8'h00;
            14'd5678: data <= 8'h00;
            14'd5679: data <= 8'h00;
            14'd5680: data <= 8'h00;
            14'd5681: data <= 8'h00;
            14'd5682: data <= 8'h00;
            14'd5683: data <= 8'h00;
            14'd5684: data <= 8'h00;
            14'd5685: data <= 8'h00;
            14'd5686: data <= 8'h0F;
            14'd5687: data <= 8'hFF;
            14'd5688: data <= 8'hFF;
            14'd5689: data <= 8'hFF;
            14'd5690: data <= 8'hFF;
            14'd5691: data <= 8'hFF;
            14'd5692: data <= 8'hFF;
            14'd5693: data <= 8'hFF;
            14'd5694: data <= 8'hFF;
            14'd5695: data <= 8'hFF;
            14'd5696: data <= 8'hFF;
            14'd5697: data <= 8'hFF;
            14'd5698: data <= 8'hFF;
            14'd5699: data <= 8'hFC;
            14'd5700: data <= 8'h3F;
            14'd5701: data <= 8'h0F;
            14'd5702: data <= 8'hF8;
            14'd5703: data <= 8'h3F;
            14'd5704: data <= 8'hFF;
            14'd5705: data <= 8'hFF;
            14'd5706: data <= 8'hFF;
            14'd5707: data <= 8'hFF;
            14'd5708: data <= 8'hFF;
            14'd5709: data <= 8'hFF;
            14'd5710: data <= 8'hFF;
            14'd5711: data <= 8'hFF;
            14'd5712: data <= 8'hFF;
            14'd5713: data <= 8'hF0;
            14'd5714: data <= 8'h00;
            14'd5715: data <= 8'h00;
            14'd5716: data <= 8'h00;
            14'd5717: data <= 8'h00;
            14'd5718: data <= 8'h00;
            14'd5719: data <= 8'h00;
            14'd5720: data <= 8'h00;
            14'd5721: data <= 8'h00;
            14'd5722: data <= 8'h00;
            14'd5723: data <= 8'h00;
            14'd5724: data <= 8'h00;
            14'd5725: data <= 8'h00;
            14'd5726: data <= 8'h0F;
            14'd5727: data <= 8'hFF;
            14'd5728: data <= 8'hFF;
            14'd5729: data <= 8'hFF;
            14'd5730: data <= 8'hFF;
            14'd5731: data <= 8'hFF;
            14'd5732: data <= 8'hFF;
            14'd5733: data <= 8'hFF;
            14'd5734: data <= 8'hFF;
            14'd5735: data <= 8'hFF;
            14'd5736: data <= 8'hFF;
            14'd5737: data <= 8'hFF;
            14'd5738: data <= 8'hDF;
            14'd5739: data <= 8'hF8;
            14'd5740: data <= 8'h7E;
            14'd5741: data <= 8'h0F;
            14'd5742: data <= 8'hF0;
            14'd5743: data <= 8'h7F;
            14'd5744: data <= 8'hFF;
            14'd5745: data <= 8'hFF;
            14'd5746: data <= 8'hFF;
            14'd5747: data <= 8'hFF;
            14'd5748: data <= 8'hFF;
            14'd5749: data <= 8'hFF;
            14'd5750: data <= 8'hFF;
            14'd5751: data <= 8'hFF;
            14'd5752: data <= 8'hFF;
            14'd5753: data <= 8'hF0;
            14'd5754: data <= 8'h00;
            14'd5755: data <= 8'h00;
            14'd5756: data <= 8'h00;
            14'd5757: data <= 8'h00;
            14'd5758: data <= 8'h00;
            14'd5759: data <= 8'h00;
            14'd5760: data <= 8'h00;
            14'd5761: data <= 8'h00;
            14'd5762: data <= 8'h00;
            14'd5763: data <= 8'h00;
            14'd5764: data <= 8'h00;
            14'd5765: data <= 8'h00;
            14'd5766: data <= 8'h0F;
            14'd5767: data <= 8'hFF;
            14'd5768: data <= 8'hFF;
            14'd5769: data <= 8'hFF;
            14'd5770: data <= 8'hFF;
            14'd5771: data <= 8'hFF;
            14'd5772: data <= 8'hFF;
            14'd5773: data <= 8'hFF;
            14'd5774: data <= 8'hFF;
            14'd5775: data <= 8'hFF;
            14'd5776: data <= 8'hFF;
            14'd5777: data <= 8'hFF;
            14'd5778: data <= 8'hFF;
            14'd5779: data <= 8'hFD;
            14'd5780: data <= 8'hFE;
            14'd5781: data <= 8'h1F;
            14'd5782: data <= 8'hF0;
            14'd5783: data <= 8'hFF;
            14'd5784: data <= 8'hFF;
            14'd5785: data <= 8'hFF;
            14'd5786: data <= 8'hFF;
            14'd5787: data <= 8'hFF;
            14'd5788: data <= 8'hFF;
            14'd5789: data <= 8'hFF;
            14'd5790: data <= 8'hFF;
            14'd5791: data <= 8'hFF;
            14'd5792: data <= 8'hFF;
            14'd5793: data <= 8'hF0;
            14'd5794: data <= 8'h00;
            14'd5795: data <= 8'h00;
            14'd5796: data <= 8'h00;
            14'd5797: data <= 8'h00;
            14'd5798: data <= 8'h00;
            14'd5799: data <= 8'h00;
            14'd5800: data <= 8'h00;
            14'd5801: data <= 8'h00;
            14'd5802: data <= 8'h00;
            14'd5803: data <= 8'h00;
            14'd5804: data <= 8'h00;
            14'd5805: data <= 8'h00;
            14'd5806: data <= 8'h0F;
            14'd5807: data <= 8'hFF;
            14'd5808: data <= 8'hFF;
            14'd5809: data <= 8'hFF;
            14'd5810: data <= 8'hFF;
            14'd5811: data <= 8'hFF;
            14'd5812: data <= 8'hFF;
            14'd5813: data <= 8'hFF;
            14'd5814: data <= 8'hFF;
            14'd5815: data <= 8'hFF;
            14'd5816: data <= 8'hFF;
            14'd5817: data <= 8'hFF;
            14'd5818: data <= 8'hFF;
            14'd5819: data <= 8'hFF;
            14'd5820: data <= 8'hFC;
            14'd5821: data <= 8'h1F;
            14'd5822: data <= 8'hE1;
            14'd5823: data <= 8'hFF;
            14'd5824: data <= 8'hFF;
            14'd5825: data <= 8'hFF;
            14'd5826: data <= 8'hFF;
            14'd5827: data <= 8'hFF;
            14'd5828: data <= 8'hFF;
            14'd5829: data <= 8'hFF;
            14'd5830: data <= 8'hFF;
            14'd5831: data <= 8'hFF;
            14'd5832: data <= 8'hFF;
            14'd5833: data <= 8'hF0;
            14'd5834: data <= 8'h00;
            14'd5835: data <= 8'h00;
            14'd5836: data <= 8'h00;
            14'd5837: data <= 8'h00;
            14'd5838: data <= 8'h00;
            14'd5839: data <= 8'h00;
            14'd5840: data <= 8'h00;
            14'd5841: data <= 8'h00;
            14'd5842: data <= 8'h00;
            14'd5843: data <= 8'h00;
            14'd5844: data <= 8'h00;
            14'd5845: data <= 8'h00;
            14'd5846: data <= 8'h0F;
            14'd5847: data <= 8'hFF;
            14'd5848: data <= 8'hFF;
            14'd5849: data <= 8'hFF;
            14'd5850: data <= 8'hFF;
            14'd5851: data <= 8'hFF;
            14'd5852: data <= 8'hFF;
            14'd5853: data <= 8'hFF;
            14'd5854: data <= 8'hFF;
            14'd5855: data <= 8'hFF;
            14'd5856: data <= 8'hFF;
            14'd5857: data <= 8'hFF;
            14'd5858: data <= 8'hFF;
            14'd5859: data <= 8'hFF;
            14'd5860: data <= 8'hEC;
            14'd5861: data <= 8'h3F;
            14'd5862: data <= 8'hC1;
            14'd5863: data <= 8'hFF;
            14'd5864: data <= 8'hFF;
            14'd5865: data <= 8'hFF;
            14'd5866: data <= 8'hFF;
            14'd5867: data <= 8'hFF;
            14'd5868: data <= 8'hFF;
            14'd5869: data <= 8'hFF;
            14'd5870: data <= 8'hFF;
            14'd5871: data <= 8'hFF;
            14'd5872: data <= 8'hFF;
            14'd5873: data <= 8'hF0;
            14'd5874: data <= 8'h00;
            14'd5875: data <= 8'h00;
            14'd5876: data <= 8'h00;
            14'd5877: data <= 8'h00;
            14'd5878: data <= 8'h00;
            14'd5879: data <= 8'h00;
            14'd5880: data <= 8'h00;
            14'd5881: data <= 8'h00;
            14'd5882: data <= 8'h00;
            14'd5883: data <= 8'h00;
            14'd5884: data <= 8'h00;
            14'd5885: data <= 8'h00;
            14'd5886: data <= 8'h0F;
            14'd5887: data <= 8'hFF;
            14'd5888: data <= 8'hFF;
            14'd5889: data <= 8'hFF;
            14'd5890: data <= 8'hFF;
            14'd5891: data <= 8'hFF;
            14'd5892: data <= 8'hFF;
            14'd5893: data <= 8'hFF;
            14'd5894: data <= 8'hFF;
            14'd5895: data <= 8'hFF;
            14'd5896: data <= 8'hFF;
            14'd5897: data <= 8'hFF;
            14'd5898: data <= 8'hFF;
            14'd5899: data <= 8'hFF;
            14'd5900: data <= 8'hF8;
            14'd5901: data <= 8'h7F;
            14'd5902: data <= 8'h83;
            14'd5903: data <= 8'hFF;
            14'd5904: data <= 8'hFF;
            14'd5905: data <= 8'hFF;
            14'd5906: data <= 8'hFF;
            14'd5907: data <= 8'hFF;
            14'd5908: data <= 8'hFF;
            14'd5909: data <= 8'hFF;
            14'd5910: data <= 8'hFF;
            14'd5911: data <= 8'hFF;
            14'd5912: data <= 8'hFF;
            14'd5913: data <= 8'hF0;
            14'd5914: data <= 8'h00;
            14'd5915: data <= 8'h00;
            14'd5916: data <= 8'h00;
            14'd5917: data <= 8'h00;
            14'd5918: data <= 8'h00;
            14'd5919: data <= 8'h00;
            14'd5920: data <= 8'h00;
            14'd5921: data <= 8'h00;
            14'd5922: data <= 8'h00;
            14'd5923: data <= 8'h00;
            14'd5924: data <= 8'h00;
            14'd5925: data <= 8'h00;
            14'd5926: data <= 8'h0F;
            14'd5927: data <= 8'hFF;
            14'd5928: data <= 8'hFF;
            14'd5929: data <= 8'hFF;
            14'd5930: data <= 8'hFF;
            14'd5931: data <= 8'hFF;
            14'd5932: data <= 8'hFF;
            14'd5933: data <= 8'hFF;
            14'd5934: data <= 8'hFF;
            14'd5935: data <= 8'hFF;
            14'd5936: data <= 8'hFF;
            14'd5937: data <= 8'hFF;
            14'd5938: data <= 8'hFF;
            14'd5939: data <= 8'hFF;
            14'd5940: data <= 8'hF8;
            14'd5941: data <= 8'hFF;
            14'd5942: data <= 8'h87;
            14'd5943: data <= 8'hFF;
            14'd5944: data <= 8'hFF;
            14'd5945: data <= 8'hFF;
            14'd5946: data <= 8'hFF;
            14'd5947: data <= 8'hFF;
            14'd5948: data <= 8'hFF;
            14'd5949: data <= 8'hFF;
            14'd5950: data <= 8'hFF;
            14'd5951: data <= 8'hFF;
            14'd5952: data <= 8'hFF;
            14'd5953: data <= 8'hF0;
            14'd5954: data <= 8'h00;
            14'd5955: data <= 8'h00;
            14'd5956: data <= 8'h00;
            14'd5957: data <= 8'h00;
            14'd5958: data <= 8'h00;
            14'd5959: data <= 8'h00;
            14'd5960: data <= 8'h00;
            14'd5961: data <= 8'h00;
            14'd5962: data <= 8'h00;
            14'd5963: data <= 8'h00;
            14'd5964: data <= 8'h00;
            14'd5965: data <= 8'h00;
            14'd5966: data <= 8'h0F;
            14'd5967: data <= 8'hFF;
            14'd5968: data <= 8'hFF;
            14'd5969: data <= 8'hFF;
            14'd5970: data <= 8'hFF;
            14'd5971: data <= 8'hFF;
            14'd5972: data <= 8'hFF;
            14'd5973: data <= 8'hFF;
            14'd5974: data <= 8'hFF;
            14'd5975: data <= 8'hFF;
            14'd5976: data <= 8'hFF;
            14'd5977: data <= 8'hFF;
            14'd5978: data <= 8'hFF;
            14'd5979: data <= 8'hFF;
            14'd5980: data <= 8'hF1;
            14'd5981: data <= 8'hFF;
            14'd5982: data <= 8'h07;
            14'd5983: data <= 8'hFF;
            14'd5984: data <= 8'hFF;
            14'd5985: data <= 8'hFF;
            14'd5986: data <= 8'hFF;
            14'd5987: data <= 8'hFF;
            14'd5988: data <= 8'hFF;
            14'd5989: data <= 8'hFF;
            14'd5990: data <= 8'hFF;
            14'd5991: data <= 8'hFF;
            14'd5992: data <= 8'hFF;
            14'd5993: data <= 8'hF0;
            14'd5994: data <= 8'h00;
            14'd5995: data <= 8'h00;
            14'd5996: data <= 8'h00;
            14'd5997: data <= 8'h00;
            14'd5998: data <= 8'h00;
            14'd5999: data <= 8'h00;
            14'd6000: data <= 8'h00;
            14'd6001: data <= 8'h00;
            14'd6002: data <= 8'h00;
            14'd6003: data <= 8'h00;
            14'd6004: data <= 8'h00;
            14'd6005: data <= 8'h00;
            14'd6006: data <= 8'h0F;
            14'd6007: data <= 8'hFF;
            14'd6008: data <= 8'hFF;
            14'd6009: data <= 8'hFF;
            14'd6010: data <= 8'hFF;
            14'd6011: data <= 8'hFF;
            14'd6012: data <= 8'hFF;
            14'd6013: data <= 8'hFF;
            14'd6014: data <= 8'hFF;
            14'd6015: data <= 8'hFF;
            14'd6016: data <= 8'hFF;
            14'd6017: data <= 8'hFF;
            14'd6018: data <= 8'h0F;
            14'd6019: data <= 8'hFF;
            14'd6020: data <= 8'hF3;
            14'd6021: data <= 8'hFE;
            14'd6022: data <= 8'h0F;
            14'd6023: data <= 8'hFF;
            14'd6024: data <= 8'hFF;
            14'd6025: data <= 8'hFF;
            14'd6026: data <= 8'hFF;
            14'd6027: data <= 8'hFF;
            14'd6028: data <= 8'hFF;
            14'd6029: data <= 8'hFF;
            14'd6030: data <= 8'hFF;
            14'd6031: data <= 8'hFF;
            14'd6032: data <= 8'hFF;
            14'd6033: data <= 8'hF0;
            14'd6034: data <= 8'h00;
            14'd6035: data <= 8'h00;
            14'd6036: data <= 8'h00;
            14'd6037: data <= 8'h00;
            14'd6038: data <= 8'h00;
            14'd6039: data <= 8'h00;
            14'd6040: data <= 8'h00;
            14'd6041: data <= 8'h00;
            14'd6042: data <= 8'h00;
            14'd6043: data <= 8'h00;
            14'd6044: data <= 8'h00;
            14'd6045: data <= 8'h00;
            14'd6046: data <= 8'h0F;
            14'd6047: data <= 8'hFF;
            14'd6048: data <= 8'hFF;
            14'd6049: data <= 8'hFF;
            14'd6050: data <= 8'hFF;
            14'd6051: data <= 8'hFF;
            14'd6052: data <= 8'hFF;
            14'd6053: data <= 8'hFF;
            14'd6054: data <= 8'hFF;
            14'd6055: data <= 8'hFF;
            14'd6056: data <= 8'hFF;
            14'd6057: data <= 8'hF8;
            14'd6058: data <= 8'h03;
            14'd6059: data <= 8'hFF;
            14'd6060: data <= 8'hF7;
            14'd6061: data <= 8'hFE;
            14'd6062: data <= 8'h1F;
            14'd6063: data <= 8'hFF;
            14'd6064: data <= 8'hFF;
            14'd6065: data <= 8'hFF;
            14'd6066: data <= 8'hFF;
            14'd6067: data <= 8'hFF;
            14'd6068: data <= 8'hFF;
            14'd6069: data <= 8'hFF;
            14'd6070: data <= 8'hFF;
            14'd6071: data <= 8'hFF;
            14'd6072: data <= 8'hFF;
            14'd6073: data <= 8'hF0;
            14'd6074: data <= 8'h00;
            14'd6075: data <= 8'h00;
            14'd6076: data <= 8'h00;
            14'd6077: data <= 8'h00;
            14'd6078: data <= 8'h00;
            14'd6079: data <= 8'h00;
            14'd6080: data <= 8'h00;
            14'd6081: data <= 8'h00;
            14'd6082: data <= 8'h00;
            14'd6083: data <= 8'h00;
            14'd6084: data <= 8'h00;
            14'd6085: data <= 8'h00;
            14'd6086: data <= 8'h0F;
            14'd6087: data <= 8'hFF;
            14'd6088: data <= 8'hFF;
            14'd6089: data <= 8'hFF;
            14'd6090: data <= 8'hFF;
            14'd6091: data <= 8'hFF;
            14'd6092: data <= 8'hFF;
            14'd6093: data <= 8'hFF;
            14'd6094: data <= 8'hFF;
            14'd6095: data <= 8'hFF;
            14'd6096: data <= 8'hF1;
            14'd6097: data <= 8'hF0;
            14'd6098: data <= 8'h01;
            14'd6099: data <= 8'hFF;
            14'd6100: data <= 8'hFF;
            14'd6101: data <= 8'hFC;
            14'd6102: data <= 8'h1F;
            14'd6103: data <= 8'hFF;
            14'd6104: data <= 8'hFF;
            14'd6105: data <= 8'hFF;
            14'd6106: data <= 8'hFF;
            14'd6107: data <= 8'hFF;
            14'd6108: data <= 8'hFF;
            14'd6109: data <= 8'hFF;
            14'd6110: data <= 8'hFF;
            14'd6111: data <= 8'hFF;
            14'd6112: data <= 8'hFF;
            14'd6113: data <= 8'hF0;
            14'd6114: data <= 8'h00;
            14'd6115: data <= 8'h00;
            14'd6116: data <= 8'h00;
            14'd6117: data <= 8'h00;
            14'd6118: data <= 8'h00;
            14'd6119: data <= 8'h00;
            14'd6120: data <= 8'h00;
            14'd6121: data <= 8'h00;
            14'd6122: data <= 8'h00;
            14'd6123: data <= 8'h00;
            14'd6124: data <= 8'h00;
            14'd6125: data <= 8'h00;
            14'd6126: data <= 8'h0F;
            14'd6127: data <= 8'hFF;
            14'd6128: data <= 8'hFF;
            14'd6129: data <= 8'hFF;
            14'd6130: data <= 8'hFF;
            14'd6131: data <= 8'hFF;
            14'd6132: data <= 8'hFF;
            14'd6133: data <= 8'hFF;
            14'd6134: data <= 8'hFF;
            14'd6135: data <= 8'hFF;
            14'd6136: data <= 8'hC0;
            14'd6137: data <= 8'h30;
            14'd6138: data <= 8'h01;
            14'd6139: data <= 8'hFF;
            14'd6140: data <= 8'hFF;
            14'd6141: data <= 8'hF8;
            14'd6142: data <= 8'h3F;
            14'd6143: data <= 8'hFF;
            14'd6144: data <= 8'hFF;
            14'd6145: data <= 8'hFF;
            14'd6146: data <= 8'hFF;
            14'd6147: data <= 8'hFF;
            14'd6148: data <= 8'hFF;
            14'd6149: data <= 8'hFF;
            14'd6150: data <= 8'hFF;
            14'd6151: data <= 8'hFF;
            14'd6152: data <= 8'hFF;
            14'd6153: data <= 8'hF0;
            14'd6154: data <= 8'h00;
            14'd6155: data <= 8'h00;
            14'd6156: data <= 8'h00;
            14'd6157: data <= 8'h00;
            14'd6158: data <= 8'h00;
            14'd6159: data <= 8'h00;
            14'd6160: data <= 8'h00;
            14'd6161: data <= 8'h00;
            14'd6162: data <= 8'h00;
            14'd6163: data <= 8'h00;
            14'd6164: data <= 8'h00;
            14'd6165: data <= 8'h00;
            14'd6166: data <= 8'h0F;
            14'd6167: data <= 8'hFF;
            14'd6168: data <= 8'hFF;
            14'd6169: data <= 8'hFF;
            14'd6170: data <= 8'hFF;
            14'd6171: data <= 8'hFF;
            14'd6172: data <= 8'hFF;
            14'd6173: data <= 8'hFF;
            14'd6174: data <= 8'hFF;
            14'd6175: data <= 8'hFF;
            14'd6176: data <= 8'h00;
            14'd6177: data <= 8'h00;
            14'd6178: data <= 8'h00;
            14'd6179: data <= 8'hFF;
            14'd6180: data <= 8'hFF;
            14'd6181: data <= 8'hF8;
            14'd6182: data <= 8'h7F;
            14'd6183: data <= 8'hFF;
            14'd6184: data <= 8'hFF;
            14'd6185: data <= 8'hFF;
            14'd6186: data <= 8'hFF;
            14'd6187: data <= 8'hFF;
            14'd6188: data <= 8'hFF;
            14'd6189: data <= 8'hFF;
            14'd6190: data <= 8'hFF;
            14'd6191: data <= 8'hFF;
            14'd6192: data <= 8'hFF;
            14'd6193: data <= 8'hF0;
            14'd6194: data <= 8'h00;
            14'd6195: data <= 8'h00;
            14'd6196: data <= 8'h00;
            14'd6197: data <= 8'h00;
            14'd6198: data <= 8'h00;
            14'd6199: data <= 8'h00;
            14'd6200: data <= 8'h00;
            14'd6201: data <= 8'h00;
            14'd6202: data <= 8'h00;
            14'd6203: data <= 8'h00;
            14'd6204: data <= 8'h00;
            14'd6205: data <= 8'h00;
            14'd6206: data <= 8'h0F;
            14'd6207: data <= 8'hFF;
            14'd6208: data <= 8'hFF;
            14'd6209: data <= 8'hFF;
            14'd6210: data <= 8'hFF;
            14'd6211: data <= 8'hFF;
            14'd6212: data <= 8'hFF;
            14'd6213: data <= 8'hFF;
            14'd6214: data <= 8'hFF;
            14'd6215: data <= 8'hFF;
            14'd6216: data <= 8'h00;
            14'd6217: data <= 8'h00;
            14'd6218: data <= 8'h60;
            14'd6219: data <= 8'hFF;
            14'd6220: data <= 8'hFF;
            14'd6221: data <= 8'hF0;
            14'd6222: data <= 8'hFF;
            14'd6223: data <= 8'hFF;
            14'd6224: data <= 8'hFF;
            14'd6225: data <= 8'hFF;
            14'd6226: data <= 8'hFF;
            14'd6227: data <= 8'hFF;
            14'd6228: data <= 8'hFF;
            14'd6229: data <= 8'hFF;
            14'd6230: data <= 8'hFF;
            14'd6231: data <= 8'hFF;
            14'd6232: data <= 8'hFF;
            14'd6233: data <= 8'hF0;
            14'd6234: data <= 8'h00;
            14'd6235: data <= 8'h00;
            14'd6236: data <= 8'h00;
            14'd6237: data <= 8'h00;
            14'd6238: data <= 8'h00;
            14'd6239: data <= 8'h00;
            14'd6240: data <= 8'h00;
            14'd6241: data <= 8'h00;
            14'd6242: data <= 8'h00;
            14'd6243: data <= 8'h00;
            14'd6244: data <= 8'h00;
            14'd6245: data <= 8'h00;
            14'd6246: data <= 8'h0F;
            14'd6247: data <= 8'hFF;
            14'd6248: data <= 8'hFF;
            14'd6249: data <= 8'hFF;
            14'd6250: data <= 8'hFF;
            14'd6251: data <= 8'hFF;
            14'd6252: data <= 8'hFF;
            14'd6253: data <= 8'hFF;
            14'd6254: data <= 8'hFF;
            14'd6255: data <= 8'hFE;
            14'd6256: data <= 8'h06;
            14'd6257: data <= 8'h01;
            14'd6258: data <= 8'hF0;
            14'd6259: data <= 8'hFF;
            14'd6260: data <= 8'hFF;
            14'd6261: data <= 8'hF1;
            14'd6262: data <= 8'hFF;
            14'd6263: data <= 8'hFF;
            14'd6264: data <= 8'hFF;
            14'd6265: data <= 8'hFF;
            14'd6266: data <= 8'hFF;
            14'd6267: data <= 8'hFF;
            14'd6268: data <= 8'hFF;
            14'd6269: data <= 8'hFF;
            14'd6270: data <= 8'hFF;
            14'd6271: data <= 8'hFF;
            14'd6272: data <= 8'hFF;
            14'd6273: data <= 8'hF0;
            14'd6274: data <= 8'h00;
            14'd6275: data <= 8'h00;
            14'd6276: data <= 8'h00;
            14'd6277: data <= 8'h00;
            14'd6278: data <= 8'h00;
            14'd6279: data <= 8'h00;
            14'd6280: data <= 8'h00;
            14'd6281: data <= 8'h00;
            14'd6282: data <= 8'h00;
            14'd6283: data <= 8'h00;
            14'd6284: data <= 8'h00;
            14'd6285: data <= 8'h00;
            14'd6286: data <= 8'h0F;
            14'd6287: data <= 8'hFF;
            14'd6288: data <= 8'hFF;
            14'd6289: data <= 8'hFF;
            14'd6290: data <= 8'hFF;
            14'd6291: data <= 8'hFF;
            14'd6292: data <= 8'hFF;
            14'd6293: data <= 8'hFF;
            14'd6294: data <= 8'hFF;
            14'd6295: data <= 8'hFE;
            14'd6296: data <= 8'h0F;
            14'd6297: data <= 8'h83;
            14'd6298: data <= 8'hF0;
            14'd6299: data <= 8'hFF;
            14'd6300: data <= 8'hFF;
            14'd6301: data <= 8'hE3;
            14'd6302: data <= 8'hFF;
            14'd6303: data <= 8'hFF;
            14'd6304: data <= 8'hFF;
            14'd6305: data <= 8'hFF;
            14'd6306: data <= 8'hFF;
            14'd6307: data <= 8'hFF;
            14'd6308: data <= 8'hFF;
            14'd6309: data <= 8'hFF;
            14'd6310: data <= 8'hFF;
            14'd6311: data <= 8'hFF;
            14'd6312: data <= 8'hFF;
            14'd6313: data <= 8'hF0;
            14'd6314: data <= 8'h00;
            14'd6315: data <= 8'h00;
            14'd6316: data <= 8'h00;
            14'd6317: data <= 8'h00;
            14'd6318: data <= 8'h00;
            14'd6319: data <= 8'h00;
            14'd6320: data <= 8'h00;
            14'd6321: data <= 8'h00;
            14'd6322: data <= 8'h00;
            14'd6323: data <= 8'h00;
            14'd6324: data <= 8'h00;
            14'd6325: data <= 8'h00;
            14'd6326: data <= 8'h0F;
            14'd6327: data <= 8'hFF;
            14'd6328: data <= 8'hFF;
            14'd6329: data <= 8'hFF;
            14'd6330: data <= 8'hFF;
            14'd6331: data <= 8'hFF;
            14'd6332: data <= 8'hFF;
            14'd6333: data <= 8'hFF;
            14'd6334: data <= 8'hFF;
            14'd6335: data <= 8'hFE;
            14'd6336: data <= 8'h0F;
            14'd6337: data <= 8'hE7;
            14'd6338: data <= 8'hF0;
            14'd6339: data <= 8'hFF;
            14'd6340: data <= 8'hFF;
            14'd6341: data <= 8'hE3;
            14'd6342: data <= 8'hFF;
            14'd6343: data <= 8'hFF;
            14'd6344: data <= 8'hFF;
            14'd6345: data <= 8'hFF;
            14'd6346: data <= 8'hFF;
            14'd6347: data <= 8'hFF;
            14'd6348: data <= 8'hFF;
            14'd6349: data <= 8'hFF;
            14'd6350: data <= 8'hFF;
            14'd6351: data <= 8'hFF;
            14'd6352: data <= 8'hFF;
            14'd6353: data <= 8'hF0;
            14'd6354: data <= 8'h00;
            14'd6355: data <= 8'h00;
            14'd6356: data <= 8'h00;
            14'd6357: data <= 8'h00;
            14'd6358: data <= 8'h00;
            14'd6359: data <= 8'h00;
            14'd6360: data <= 8'h00;
            14'd6361: data <= 8'h00;
            14'd6362: data <= 8'h00;
            14'd6363: data <= 8'h00;
            14'd6364: data <= 8'h00;
            14'd6365: data <= 8'h00;
            14'd6366: data <= 8'h0F;
            14'd6367: data <= 8'hFF;
            14'd6368: data <= 8'hFF;
            14'd6369: data <= 8'hFF;
            14'd6370: data <= 8'hFF;
            14'd6371: data <= 8'hFF;
            14'd6372: data <= 8'hFF;
            14'd6373: data <= 8'hFF;
            14'd6374: data <= 8'hFF;
            14'd6375: data <= 8'hFC;
            14'd6376: data <= 8'h1F;
            14'd6377: data <= 8'hBF;
            14'd6378: data <= 8'hE0;
            14'd6379: data <= 8'hFF;
            14'd6380: data <= 8'hFF;
            14'd6381: data <= 8'hC7;
            14'd6382: data <= 8'hFF;
            14'd6383: data <= 8'hFF;
            14'd6384: data <= 8'hFF;
            14'd6385: data <= 8'hFF;
            14'd6386: data <= 8'hFF;
            14'd6387: data <= 8'hFF;
            14'd6388: data <= 8'hFF;
            14'd6389: data <= 8'hFF;
            14'd6390: data <= 8'hFF;
            14'd6391: data <= 8'hFF;
            14'd6392: data <= 8'hFF;
            14'd6393: data <= 8'hF0;
            14'd6394: data <= 8'h00;
            14'd6395: data <= 8'h00;
            14'd6396: data <= 8'h00;
            14'd6397: data <= 8'h00;
            14'd6398: data <= 8'h00;
            14'd6399: data <= 8'h00;
            14'd6400: data <= 8'h00;
            14'd6401: data <= 8'h00;
            14'd6402: data <= 8'h00;
            14'd6403: data <= 8'h00;
            14'd6404: data <= 8'h00;
            14'd6405: data <= 8'h00;
            14'd6406: data <= 8'h0F;
            14'd6407: data <= 8'hFF;
            14'd6408: data <= 8'hFF;
            14'd6409: data <= 8'hFF;
            14'd6410: data <= 8'hFF;
            14'd6411: data <= 8'hFF;
            14'd6412: data <= 8'hFF;
            14'd6413: data <= 8'hFF;
            14'd6414: data <= 8'hFF;
            14'd6415: data <= 8'hFE;
            14'd6416: data <= 8'h0F;
            14'd6417: data <= 8'hFF;
            14'd6418: data <= 8'hE0;
            14'd6419: data <= 8'hFF;
            14'd6420: data <= 8'hFF;
            14'd6421: data <= 8'h8F;
            14'd6422: data <= 8'hFF;
            14'd6423: data <= 8'hFF;
            14'd6424: data <= 8'hFF;
            14'd6425: data <= 8'hFF;
            14'd6426: data <= 8'hFF;
            14'd6427: data <= 8'hFF;
            14'd6428: data <= 8'hFF;
            14'd6429: data <= 8'hFF;
            14'd6430: data <= 8'hFF;
            14'd6431: data <= 8'hFF;
            14'd6432: data <= 8'hFF;
            14'd6433: data <= 8'hF0;
            14'd6434: data <= 8'h00;
            14'd6435: data <= 8'h00;
            14'd6436: data <= 8'h00;
            14'd6437: data <= 8'h00;
            14'd6438: data <= 8'h00;
            14'd6439: data <= 8'h00;
            14'd6440: data <= 8'h00;
            14'd6441: data <= 8'h00;
            14'd6442: data <= 8'h00;
            14'd6443: data <= 8'h00;
            14'd6444: data <= 8'h00;
            14'd6445: data <= 8'h00;
            14'd6446: data <= 8'h0F;
            14'd6447: data <= 8'hFF;
            14'd6448: data <= 8'hFF;
            14'd6449: data <= 8'hFF;
            14'd6450: data <= 8'hFF;
            14'd6451: data <= 8'hFF;
            14'd6452: data <= 8'hFF;
            14'd6453: data <= 8'hFF;
            14'd6454: data <= 8'hFF;
            14'd6455: data <= 8'hFE;
            14'd6456: data <= 8'h07;
            14'd6457: data <= 8'hFF;
            14'd6458: data <= 8'hE0;
            14'd6459: data <= 8'hFF;
            14'd6460: data <= 8'hFF;
            14'd6461: data <= 8'h9F;
            14'd6462: data <= 8'hFF;
            14'd6463: data <= 8'hFF;
            14'd6464: data <= 8'hFF;
            14'd6465: data <= 8'hFF;
            14'd6466: data <= 8'hFF;
            14'd6467: data <= 8'hFF;
            14'd6468: data <= 8'hFF;
            14'd6469: data <= 8'hFF;
            14'd6470: data <= 8'hFF;
            14'd6471: data <= 8'hFF;
            14'd6472: data <= 8'hFF;
            14'd6473: data <= 8'hF0;
            14'd6474: data <= 8'h00;
            14'd6475: data <= 8'h00;
            14'd6476: data <= 8'h00;
            14'd6477: data <= 8'h00;
            14'd6478: data <= 8'h00;
            14'd6479: data <= 8'h00;
            14'd6480: data <= 8'h00;
            14'd6481: data <= 8'h00;
            14'd6482: data <= 8'h00;
            14'd6483: data <= 8'h00;
            14'd6484: data <= 8'h00;
            14'd6485: data <= 8'h00;
            14'd6486: data <= 8'h0F;
            14'd6487: data <= 8'hFF;
            14'd6488: data <= 8'hFF;
            14'd6489: data <= 8'hFF;
            14'd6490: data <= 8'hFF;
            14'd6491: data <= 8'hFF;
            14'd6492: data <= 8'hFF;
            14'd6493: data <= 8'hFF;
            14'd6494: data <= 8'hFF;
            14'd6495: data <= 8'hFE;
            14'd6496: data <= 8'h07;
            14'd6497: data <= 8'hFF;
            14'd6498: data <= 8'hC1;
            14'd6499: data <= 8'hFF;
            14'd6500: data <= 8'hFF;
            14'd6501: data <= 8'h3F;
            14'd6502: data <= 8'hFF;
            14'd6503: data <= 8'hFF;
            14'd6504: data <= 8'hFF;
            14'd6505: data <= 8'hFF;
            14'd6506: data <= 8'hFF;
            14'd6507: data <= 8'hFF;
            14'd6508: data <= 8'hFF;
            14'd6509: data <= 8'hFF;
            14'd6510: data <= 8'hFF;
            14'd6511: data <= 8'hFF;
            14'd6512: data <= 8'hFF;
            14'd6513: data <= 8'hF0;
            14'd6514: data <= 8'h00;
            14'd6515: data <= 8'h00;
            14'd6516: data <= 8'h00;
            14'd6517: data <= 8'h00;
            14'd6518: data <= 8'h00;
            14'd6519: data <= 8'h00;
            14'd6520: data <= 8'h00;
            14'd6521: data <= 8'h00;
            14'd6522: data <= 8'h00;
            14'd6523: data <= 8'h00;
            14'd6524: data <= 8'h00;
            14'd6525: data <= 8'h00;
            14'd6526: data <= 8'h0F;
            14'd6527: data <= 8'hFF;
            14'd6528: data <= 8'hFF;
            14'd6529: data <= 8'hFF;
            14'd6530: data <= 8'hFF;
            14'd6531: data <= 8'hFF;
            14'd6532: data <= 8'hFF;
            14'd6533: data <= 8'hFB;
            14'd6534: data <= 8'hFF;
            14'd6535: data <= 8'hFF;
            14'd6536: data <= 8'h03;
            14'd6537: data <= 8'hFF;
            14'd6538: data <= 8'hC1;
            14'd6539: data <= 8'hFF;
            14'd6540: data <= 8'hFF;
            14'd6541: data <= 8'h3F;
            14'd6542: data <= 8'hFF;
            14'd6543: data <= 8'hFF;
            14'd6544: data <= 8'hFF;
            14'd6545: data <= 8'hFF;
            14'd6546: data <= 8'hFF;
            14'd6547: data <= 8'hFF;
            14'd6548: data <= 8'hFF;
            14'd6549: data <= 8'hFF;
            14'd6550: data <= 8'hFF;
            14'd6551: data <= 8'hFF;
            14'd6552: data <= 8'hFF;
            14'd6553: data <= 8'hF0;
            14'd6554: data <= 8'h00;
            14'd6555: data <= 8'h00;
            14'd6556: data <= 8'h00;
            14'd6557: data <= 8'h00;
            14'd6558: data <= 8'h00;
            14'd6559: data <= 8'h00;
            14'd6560: data <= 8'h00;
            14'd6561: data <= 8'h00;
            14'd6562: data <= 8'h00;
            14'd6563: data <= 8'h00;
            14'd6564: data <= 8'h00;
            14'd6565: data <= 8'h00;
            14'd6566: data <= 8'h0F;
            14'd6567: data <= 8'hFF;
            14'd6568: data <= 8'hFF;
            14'd6569: data <= 8'hFF;
            14'd6570: data <= 8'hFF;
            14'd6571: data <= 8'hFF;
            14'd6572: data <= 8'hFF;
            14'd6573: data <= 8'hFF;
            14'd6574: data <= 8'hFF;
            14'd6575: data <= 8'hFF;
            14'd6576: data <= 8'h81;
            14'd6577: data <= 8'hFF;
            14'd6578: data <= 8'h81;
            14'd6579: data <= 8'hFF;
            14'd6580: data <= 8'hFE;
            14'd6581: data <= 8'h7F;
            14'd6582: data <= 8'hFF;
            14'd6583: data <= 8'hFF;
            14'd6584: data <= 8'hFF;
            14'd6585: data <= 8'hFF;
            14'd6586: data <= 8'hFF;
            14'd6587: data <= 8'hFF;
            14'd6588: data <= 8'hFF;
            14'd6589: data <= 8'hFF;
            14'd6590: data <= 8'hFF;
            14'd6591: data <= 8'hFF;
            14'd6592: data <= 8'hFF;
            14'd6593: data <= 8'hF0;
            14'd6594: data <= 8'h00;
            14'd6595: data <= 8'h00;
            14'd6596: data <= 8'h00;
            14'd6597: data <= 8'h00;
            14'd6598: data <= 8'h00;
            14'd6599: data <= 8'h00;
            14'd6600: data <= 8'h00;
            14'd6601: data <= 8'h00;
            14'd6602: data <= 8'h00;
            14'd6603: data <= 8'h00;
            14'd6604: data <= 8'h00;
            14'd6605: data <= 8'h00;
            14'd6606: data <= 8'h0F;
            14'd6607: data <= 8'hFF;
            14'd6608: data <= 8'hFF;
            14'd6609: data <= 8'hFF;
            14'd6610: data <= 8'hFF;
            14'd6611: data <= 8'hFF;
            14'd6612: data <= 8'hFF;
            14'd6613: data <= 8'hFF;
            14'd6614: data <= 8'hFF;
            14'd6615: data <= 8'hFF;
            14'd6616: data <= 8'h80;
            14'd6617: data <= 8'hFF;
            14'd6618: data <= 8'h03;
            14'd6619: data <= 8'hFF;
            14'd6620: data <= 8'hFF;
            14'd6621: data <= 8'hFF;
            14'd6622: data <= 8'hFF;
            14'd6623: data <= 8'hFF;
            14'd6624: data <= 8'hFF;
            14'd6625: data <= 8'hFF;
            14'd6626: data <= 8'hFF;
            14'd6627: data <= 8'hFF;
            14'd6628: data <= 8'hFF;
            14'd6629: data <= 8'hFF;
            14'd6630: data <= 8'hFF;
            14'd6631: data <= 8'hFF;
            14'd6632: data <= 8'hFF;
            14'd6633: data <= 8'hF0;
            14'd6634: data <= 8'h00;
            14'd6635: data <= 8'h00;
            14'd6636: data <= 8'h00;
            14'd6637: data <= 8'h00;
            14'd6638: data <= 8'h00;
            14'd6639: data <= 8'h00;
            14'd6640: data <= 8'h00;
            14'd6641: data <= 8'h00;
            14'd6642: data <= 8'h00;
            14'd6643: data <= 8'h00;
            14'd6644: data <= 8'h00;
            14'd6645: data <= 8'h00;
            14'd6646: data <= 8'h0F;
            14'd6647: data <= 8'hBF;
            14'd6648: data <= 8'hFF;
            14'd6649: data <= 8'hFF;
            14'd6650: data <= 8'hFF;
            14'd6651: data <= 8'hFF;
            14'd6652: data <= 8'hFF;
            14'd6653: data <= 8'hFF;
            14'd6654: data <= 8'hFF;
            14'd6655: data <= 8'hFF;
            14'd6656: data <= 8'hC0;
            14'd6657: data <= 8'h7E;
            14'd6658: data <= 8'h07;
            14'd6659: data <= 8'hFF;
            14'd6660: data <= 8'hFF;
            14'd6661: data <= 8'hFF;
            14'd6662: data <= 8'hFF;
            14'd6663: data <= 8'hFF;
            14'd6664: data <= 8'hFF;
            14'd6665: data <= 8'hFF;
            14'd6666: data <= 8'hFF;
            14'd6667: data <= 8'hFF;
            14'd6668: data <= 8'hFF;
            14'd6669: data <= 8'hFF;
            14'd6670: data <= 8'hFF;
            14'd6671: data <= 8'hFF;
            14'd6672: data <= 8'hFF;
            14'd6673: data <= 8'hF0;
            14'd6674: data <= 8'h00;
            14'd6675: data <= 8'h00;
            14'd6676: data <= 8'h00;
            14'd6677: data <= 8'h00;
            14'd6678: data <= 8'h00;
            14'd6679: data <= 8'h00;
            14'd6680: data <= 8'h00;
            14'd6681: data <= 8'h00;
            14'd6682: data <= 8'h00;
            14'd6683: data <= 8'h00;
            14'd6684: data <= 8'h00;
            14'd6685: data <= 8'h00;
            14'd6686: data <= 8'h0F;
            14'd6687: data <= 8'hBF;
            14'd6688: data <= 8'hFF;
            14'd6689: data <= 8'hFF;
            14'd6690: data <= 8'hFF;
            14'd6691: data <= 8'hFF;
            14'd6692: data <= 8'hFF;
            14'd6693: data <= 8'hFF;
            14'd6694: data <= 8'hFF;
            14'd6695: data <= 8'hFF;
            14'd6696: data <= 8'hE0;
            14'd6697: data <= 8'h3C;
            14'd6698: data <= 8'h07;
            14'd6699: data <= 8'hFF;
            14'd6700: data <= 8'hFF;
            14'd6701: data <= 8'hFF;
            14'd6702: data <= 8'hFF;
            14'd6703: data <= 8'hFF;
            14'd6704: data <= 8'hFF;
            14'd6705: data <= 8'hFF;
            14'd6706: data <= 8'hFF;
            14'd6707: data <= 8'hFF;
            14'd6708: data <= 8'hFF;
            14'd6709: data <= 8'hFF;
            14'd6710: data <= 8'hFF;
            14'd6711: data <= 8'hFF;
            14'd6712: data <= 8'hFF;
            14'd6713: data <= 8'hF0;
            14'd6714: data <= 8'h00;
            14'd6715: data <= 8'h00;
            14'd6716: data <= 8'h00;
            14'd6717: data <= 8'h00;
            14'd6718: data <= 8'h00;
            14'd6719: data <= 8'h00;
            14'd6720: data <= 8'h00;
            14'd6721: data <= 8'h00;
            14'd6722: data <= 8'h00;
            14'd6723: data <= 8'h00;
            14'd6724: data <= 8'h00;
            14'd6725: data <= 8'h00;
            14'd6726: data <= 8'h0F;
            14'd6727: data <= 8'hFF;
            14'd6728: data <= 8'hFF;
            14'd6729: data <= 8'hFF;
            14'd6730: data <= 8'hFF;
            14'd6731: data <= 8'hFF;
            14'd6732: data <= 8'hFF;
            14'd6733: data <= 8'hFF;
            14'd6734: data <= 8'hFF;
            14'd6735: data <= 8'hFF;
            14'd6736: data <= 8'hF0;
            14'd6737: data <= 8'h08;
            14'd6738: data <= 8'h0F;
            14'd6739: data <= 8'hFF;
            14'd6740: data <= 8'hFF;
            14'd6741: data <= 8'hFF;
            14'd6742: data <= 8'hFF;
            14'd6743: data <= 8'hFF;
            14'd6744: data <= 8'hFF;
            14'd6745: data <= 8'hFF;
            14'd6746: data <= 8'hFF;
            14'd6747: data <= 8'hFF;
            14'd6748: data <= 8'hFF;
            14'd6749: data <= 8'hFF;
            14'd6750: data <= 8'hFF;
            14'd6751: data <= 8'hFF;
            14'd6752: data <= 8'hFF;
            14'd6753: data <= 8'hF0;
            14'd6754: data <= 8'h00;
            14'd6755: data <= 8'h00;
            14'd6756: data <= 8'h00;
            14'd6757: data <= 8'h00;
            14'd6758: data <= 8'h00;
            14'd6759: data <= 8'h00;
            14'd6760: data <= 8'h00;
            14'd6761: data <= 8'h00;
            14'd6762: data <= 8'h00;
            14'd6763: data <= 8'h00;
            14'd6764: data <= 8'h00;
            14'd6765: data <= 8'h00;
            14'd6766: data <= 8'h0F;
            14'd6767: data <= 8'hFF;
            14'd6768: data <= 8'hFF;
            14'd6769: data <= 8'hFF;
            14'd6770: data <= 8'hFF;
            14'd6771: data <= 8'hFF;
            14'd6772: data <= 8'hFF;
            14'd6773: data <= 8'hFF;
            14'd6774: data <= 8'hFF;
            14'd6775: data <= 8'hFF;
            14'd6776: data <= 8'hFC;
            14'd6777: data <= 8'h00;
            14'd6778: data <= 8'h1F;
            14'd6779: data <= 8'hFF;
            14'd6780: data <= 8'hFF;
            14'd6781: data <= 8'hFF;
            14'd6782: data <= 8'hFF;
            14'd6783: data <= 8'hFF;
            14'd6784: data <= 8'hFF;
            14'd6785: data <= 8'hFF;
            14'd6786: data <= 8'hFF;
            14'd6787: data <= 8'hFF;
            14'd6788: data <= 8'hFF;
            14'd6789: data <= 8'hFF;
            14'd6790: data <= 8'hFF;
            14'd6791: data <= 8'hFF;
            14'd6792: data <= 8'hFF;
            14'd6793: data <= 8'hF0;
            14'd6794: data <= 8'h00;
            14'd6795: data <= 8'h00;
            14'd6796: data <= 8'h00;
            14'd6797: data <= 8'h00;
            14'd6798: data <= 8'h00;
            14'd6799: data <= 8'h00;
            14'd6800: data <= 8'h00;
            14'd6801: data <= 8'h00;
            14'd6802: data <= 8'h00;
            14'd6803: data <= 8'h00;
            14'd6804: data <= 8'h00;
            14'd6805: data <= 8'h00;
            14'd6806: data <= 8'h0F;
            14'd6807: data <= 8'hFF;
            14'd6808: data <= 8'hFF;
            14'd6809: data <= 8'hFF;
            14'd6810: data <= 8'hFF;
            14'd6811: data <= 8'hFF;
            14'd6812: data <= 8'hFF;
            14'd6813: data <= 8'hFF;
            14'd6814: data <= 8'hFF;
            14'd6815: data <= 8'hFF;
            14'd6816: data <= 8'hFE;
            14'd6817: data <= 8'h00;
            14'd6818: data <= 8'h3F;
            14'd6819: data <= 8'hFF;
            14'd6820: data <= 8'hFF;
            14'd6821: data <= 8'hFF;
            14'd6822: data <= 8'hFF;
            14'd6823: data <= 8'hFF;
            14'd6824: data <= 8'hFF;
            14'd6825: data <= 8'hFF;
            14'd6826: data <= 8'hFF;
            14'd6827: data <= 8'hFF;
            14'd6828: data <= 8'hFF;
            14'd6829: data <= 8'hFF;
            14'd6830: data <= 8'hFF;
            14'd6831: data <= 8'hFF;
            14'd6832: data <= 8'hFF;
            14'd6833: data <= 8'hF0;
            14'd6834: data <= 8'h00;
            14'd6835: data <= 8'h00;
            14'd6836: data <= 8'h00;
            14'd6837: data <= 8'h00;
            14'd6838: data <= 8'h00;
            14'd6839: data <= 8'h00;
            14'd6840: data <= 8'h00;
            14'd6841: data <= 8'h00;
            14'd6842: data <= 8'h00;
            14'd6843: data <= 8'h00;
            14'd6844: data <= 8'h00;
            14'd6845: data <= 8'h00;
            14'd6846: data <= 8'h0F;
            14'd6847: data <= 8'hFF;
            14'd6848: data <= 8'hFF;
            14'd6849: data <= 8'hFF;
            14'd6850: data <= 8'hFF;
            14'd6851: data <= 8'hFF;
            14'd6852: data <= 8'hFF;
            14'd6853: data <= 8'hFF;
            14'd6854: data <= 8'hFF;
            14'd6855: data <= 8'hFF;
            14'd6856: data <= 8'hF3;
            14'd6857: data <= 8'h00;
            14'd6858: data <= 8'h7F;
            14'd6859: data <= 8'hFF;
            14'd6860: data <= 8'hFF;
            14'd6861: data <= 8'hFF;
            14'd6862: data <= 8'hFF;
            14'd6863: data <= 8'hFF;
            14'd6864: data <= 8'hFF;
            14'd6865: data <= 8'hFF;
            14'd6866: data <= 8'hFF;
            14'd6867: data <= 8'hFF;
            14'd6868: data <= 8'hFF;
            14'd6869: data <= 8'hFF;
            14'd6870: data <= 8'hFF;
            14'd6871: data <= 8'hFF;
            14'd6872: data <= 8'hFF;
            14'd6873: data <= 8'hF0;
            14'd6874: data <= 8'h00;
            14'd6875: data <= 8'h00;
            14'd6876: data <= 8'h00;
            14'd6877: data <= 8'h00;
            14'd6878: data <= 8'h00;
            14'd6879: data <= 8'h00;
            14'd6880: data <= 8'h00;
            14'd6881: data <= 8'h00;
            14'd6882: data <= 8'h00;
            14'd6883: data <= 8'h00;
            14'd6884: data <= 8'h00;
            14'd6885: data <= 8'h00;
            14'd6886: data <= 8'h0F;
            14'd6887: data <= 8'hFF;
            14'd6888: data <= 8'hFF;
            14'd6889: data <= 8'hFF;
            14'd6890: data <= 8'hFF;
            14'd6891: data <= 8'hFF;
            14'd6892: data <= 8'hFF;
            14'd6893: data <= 8'hFF;
            14'd6894: data <= 8'hFF;
            14'd6895: data <= 8'hFF;
            14'd6896: data <= 8'hF9;
            14'd6897: data <= 8'hC0;
            14'd6898: data <= 8'hFF;
            14'd6899: data <= 8'hFF;
            14'd6900: data <= 8'hFF;
            14'd6901: data <= 8'hFF;
            14'd6902: data <= 8'hFF;
            14'd6903: data <= 8'hFF;
            14'd6904: data <= 8'hFF;
            14'd6905: data <= 8'hFF;
            14'd6906: data <= 8'hFF;
            14'd6907: data <= 8'hFF;
            14'd6908: data <= 8'hFF;
            14'd6909: data <= 8'hFF;
            14'd6910: data <= 8'hFF;
            14'd6911: data <= 8'hFF;
            14'd6912: data <= 8'hFF;
            14'd6913: data <= 8'hF0;
            14'd6914: data <= 8'h00;
            14'd6915: data <= 8'h00;
            14'd6916: data <= 8'h00;
            14'd6917: data <= 8'h00;
            14'd6918: data <= 8'h00;
            14'd6919: data <= 8'h00;
            14'd6920: data <= 8'h00;
            14'd6921: data <= 8'h00;
            14'd6922: data <= 8'h00;
            14'd6923: data <= 8'h00;
            14'd6924: data <= 8'h00;
            14'd6925: data <= 8'h00;
            14'd6926: data <= 8'h0F;
            14'd6927: data <= 8'hFF;
            14'd6928: data <= 8'hFF;
            14'd6929: data <= 8'h7F;
            14'd6930: data <= 8'hFF;
            14'd6931: data <= 8'hFF;
            14'd6932: data <= 8'hFF;
            14'd6933: data <= 8'hFF;
            14'd6934: data <= 8'hFF;
            14'd6935: data <= 8'hFF;
            14'd6936: data <= 8'hFF;
            14'd6937: data <= 8'hF3;
            14'd6938: data <= 8'hFF;
            14'd6939: data <= 8'hFF;
            14'd6940: data <= 8'hFF;
            14'd6941: data <= 8'hFF;
            14'd6942: data <= 8'hFF;
            14'd6943: data <= 8'hFF;
            14'd6944: data <= 8'hFF;
            14'd6945: data <= 8'hFF;
            14'd6946: data <= 8'hFF;
            14'd6947: data <= 8'hFF;
            14'd6948: data <= 8'hFF;
            14'd6949: data <= 8'hFF;
            14'd6950: data <= 8'hFF;
            14'd6951: data <= 8'hFF;
            14'd6952: data <= 8'hFF;
            14'd6953: data <= 8'hF0;
            14'd6954: data <= 8'h00;
            14'd6955: data <= 8'h00;
            14'd6956: data <= 8'h00;
            14'd6957: data <= 8'h00;
            14'd6958: data <= 8'h00;
            14'd6959: data <= 8'h00;
            14'd6960: data <= 8'h00;
            14'd6961: data <= 8'h00;
            14'd6962: data <= 8'h00;
            14'd6963: data <= 8'h00;
            14'd6964: data <= 8'h00;
            14'd6965: data <= 8'h00;
            14'd6966: data <= 8'h0F;
            14'd6967: data <= 8'hFF;
            14'd6968: data <= 8'hFF;
            14'd6969: data <= 8'hFF;
            14'd6970: data <= 8'hFF;
            14'd6971: data <= 8'hFF;
            14'd6972: data <= 8'hFF;
            14'd6973: data <= 8'hFF;
            14'd6974: data <= 8'hFF;
            14'd6975: data <= 8'hFF;
            14'd6976: data <= 8'hFF;
            14'd6977: data <= 8'hBF;
            14'd6978: data <= 8'hFF;
            14'd6979: data <= 8'hFF;
            14'd6980: data <= 8'hFF;
            14'd6981: data <= 8'hFF;
            14'd6982: data <= 8'hFF;
            14'd6983: data <= 8'hFF;
            14'd6984: data <= 8'hFF;
            14'd6985: data <= 8'hFF;
            14'd6986: data <= 8'hFF;
            14'd6987: data <= 8'hFF;
            14'd6988: data <= 8'hFF;
            14'd6989: data <= 8'hFF;
            14'd6990: data <= 8'hFF;
            14'd6991: data <= 8'hFF;
            14'd6992: data <= 8'hFF;
            14'd6993: data <= 8'hF0;
            14'd6994: data <= 8'h00;
            14'd6995: data <= 8'h00;
            14'd6996: data <= 8'h00;
            14'd6997: data <= 8'h00;
            14'd6998: data <= 8'h00;
            14'd6999: data <= 8'h00;
            14'd7000: data <= 8'h00;
            14'd7001: data <= 8'h00;
            14'd7002: data <= 8'h00;
            14'd7003: data <= 8'h00;
            14'd7004: data <= 8'h00;
            14'd7005: data <= 8'h00;
            14'd7006: data <= 8'h0F;
            14'd7007: data <= 8'hFF;
            14'd7008: data <= 8'hFF;
            14'd7009: data <= 8'hFF;
            14'd7010: data <= 8'hFF;
            14'd7011: data <= 8'hFF;
            14'd7012: data <= 8'hFF;
            14'd7013: data <= 8'hFF;
            14'd7014: data <= 8'hFF;
            14'd7015: data <= 8'hFF;
            14'd7016: data <= 8'hFF;
            14'd7017: data <= 8'hFF;
            14'd7018: data <= 8'hFF;
            14'd7019: data <= 8'hFF;
            14'd7020: data <= 8'hFF;
            14'd7021: data <= 8'hFF;
            14'd7022: data <= 8'hFF;
            14'd7023: data <= 8'hFF;
            14'd7024: data <= 8'hFF;
            14'd7025: data <= 8'hFF;
            14'd7026: data <= 8'hFF;
            14'd7027: data <= 8'hFF;
            14'd7028: data <= 8'hFF;
            14'd7029: data <= 8'hFF;
            14'd7030: data <= 8'hFF;
            14'd7031: data <= 8'hFF;
            14'd7032: data <= 8'hFF;
            14'd7033: data <= 8'hF0;
            14'd7034: data <= 8'h00;
            14'd7035: data <= 8'h00;
            14'd7036: data <= 8'h00;
            14'd7037: data <= 8'h00;
            14'd7038: data <= 8'h00;
            14'd7039: data <= 8'h00;
            14'd7040: data <= 8'h00;
            14'd7041: data <= 8'h00;
            14'd7042: data <= 8'h00;
            14'd7043: data <= 8'h00;
            14'd7044: data <= 8'h00;
            14'd7045: data <= 8'h00;
            14'd7046: data <= 8'h0F;
            14'd7047: data <= 8'hFF;
            14'd7048: data <= 8'hFF;
            14'd7049: data <= 8'hFF;
            14'd7050: data <= 8'hFF;
            14'd7051: data <= 8'hFF;
            14'd7052: data <= 8'hFF;
            14'd7053: data <= 8'hFF;
            14'd7054: data <= 8'hFF;
            14'd7055: data <= 8'hFF;
            14'd7056: data <= 8'hFF;
            14'd7057: data <= 8'hFF;
            14'd7058: data <= 8'hFF;
            14'd7059: data <= 8'hFF;
            14'd7060: data <= 8'hFF;
            14'd7061: data <= 8'hFF;
            14'd7062: data <= 8'hFF;
            14'd7063: data <= 8'hFF;
            14'd7064: data <= 8'hFF;
            14'd7065: data <= 8'hFF;
            14'd7066: data <= 8'hFF;
            14'd7067: data <= 8'hFF;
            14'd7068: data <= 8'hFF;
            14'd7069: data <= 8'hFF;
            14'd7070: data <= 8'hFF;
            14'd7071: data <= 8'hFF;
            14'd7072: data <= 8'hFF;
            14'd7073: data <= 8'hF0;
            14'd7074: data <= 8'h00;
            14'd7075: data <= 8'h00;
            14'd7076: data <= 8'h00;
            14'd7077: data <= 8'h00;
            14'd7078: data <= 8'h00;
            14'd7079: data <= 8'h00;
            14'd7080: data <= 8'h00;
            14'd7081: data <= 8'h00;
            14'd7082: data <= 8'h00;
            14'd7083: data <= 8'h00;
            14'd7084: data <= 8'h00;
            14'd7085: data <= 8'h00;
            14'd7086: data <= 8'h0F;
            14'd7087: data <= 8'hFF;
            14'd7088: data <= 8'hFF;
            14'd7089: data <= 8'hFF;
            14'd7090: data <= 8'hFF;
            14'd7091: data <= 8'hFF;
            14'd7092: data <= 8'hFF;
            14'd7093: data <= 8'hFF;
            14'd7094: data <= 8'hFF;
            14'd7095: data <= 8'hFF;
            14'd7096: data <= 8'hFF;
            14'd7097: data <= 8'hFF;
            14'd7098: data <= 8'hFF;
            14'd7099: data <= 8'hFF;
            14'd7100: data <= 8'hFF;
            14'd7101: data <= 8'hFF;
            14'd7102: data <= 8'hFF;
            14'd7103: data <= 8'hFF;
            14'd7104: data <= 8'hFF;
            14'd7105: data <= 8'hFF;
            14'd7106: data <= 8'hFF;
            14'd7107: data <= 8'hFF;
            14'd7108: data <= 8'hFF;
            14'd7109: data <= 8'hFF;
            14'd7110: data <= 8'hFF;
            14'd7111: data <= 8'hFF;
            14'd7112: data <= 8'hFF;
            14'd7113: data <= 8'hF0;
            14'd7114: data <= 8'h00;
            14'd7115: data <= 8'h00;
            14'd7116: data <= 8'h00;
            14'd7117: data <= 8'h00;
            14'd7118: data <= 8'h00;
            14'd7119: data <= 8'h00;
            14'd7120: data <= 8'h00;
            14'd7121: data <= 8'h00;
            14'd7122: data <= 8'h00;
            14'd7123: data <= 8'h00;
            14'd7124: data <= 8'h00;
            14'd7125: data <= 8'h00;
            14'd7126: data <= 8'h0F;
            14'd7127: data <= 8'hFF;
            14'd7128: data <= 8'hFF;
            14'd7129: data <= 8'hFF;
            14'd7130: data <= 8'hFF;
            14'd7131: data <= 8'hFF;
            14'd7132: data <= 8'hFF;
            14'd7133: data <= 8'hFF;
            14'd7134: data <= 8'hFF;
            14'd7135: data <= 8'hFF;
            14'd7136: data <= 8'hFF;
            14'd7137: data <= 8'hFF;
            14'd7138: data <= 8'hFF;
            14'd7139: data <= 8'hFF;
            14'd7140: data <= 8'hFF;
            14'd7141: data <= 8'hFF;
            14'd7142: data <= 8'hFF;
            14'd7143: data <= 8'hFF;
            14'd7144: data <= 8'hFF;
            14'd7145: data <= 8'hFF;
            14'd7146: data <= 8'hFF;
            14'd7147: data <= 8'hFF;
            14'd7148: data <= 8'hFF;
            14'd7149: data <= 8'hFF;
            14'd7150: data <= 8'hFF;
            14'd7151: data <= 8'hFF;
            14'd7152: data <= 8'hFF;
            14'd7153: data <= 8'hF0;
            14'd7154: data <= 8'h00;
            14'd7155: data <= 8'h00;
            14'd7156: data <= 8'h00;
            14'd7157: data <= 8'h00;
            14'd7158: data <= 8'h00;
            14'd7159: data <= 8'h00;
            14'd7160: data <= 8'h00;
            14'd7161: data <= 8'h00;
            14'd7162: data <= 8'h00;
            14'd7163: data <= 8'h00;
            14'd7164: data <= 8'h00;
            14'd7165: data <= 8'h00;
            14'd7166: data <= 8'h0F;
            14'd7167: data <= 8'hFF;
            14'd7168: data <= 8'hFF;
            14'd7169: data <= 8'hFF;
            14'd7170: data <= 8'hFF;
            14'd7171: data <= 8'hFF;
            14'd7172: data <= 8'hFF;
            14'd7173: data <= 8'hFF;
            14'd7174: data <= 8'hFF;
            14'd7175: data <= 8'hFF;
            14'd7176: data <= 8'hFF;
            14'd7177: data <= 8'hFF;
            14'd7178: data <= 8'hFF;
            14'd7179: data <= 8'hFF;
            14'd7180: data <= 8'hFF;
            14'd7181: data <= 8'hFF;
            14'd7182: data <= 8'hFF;
            14'd7183: data <= 8'hFF;
            14'd7184: data <= 8'hFF;
            14'd7185: data <= 8'hFF;
            14'd7186: data <= 8'hFF;
            14'd7187: data <= 8'hFF;
            14'd7188: data <= 8'hFF;
            14'd7189: data <= 8'hFF;
            14'd7190: data <= 8'hFF;
            14'd7191: data <= 8'hFF;
            14'd7192: data <= 8'hFF;
            14'd7193: data <= 8'hF0;
            14'd7194: data <= 8'h00;
            14'd7195: data <= 8'h00;
            14'd7196: data <= 8'h00;
            14'd7197: data <= 8'h00;
            14'd7198: data <= 8'h00;
            14'd7199: data <= 8'h00;
            14'd7200: data <= 8'h00;
            14'd7201: data <= 8'h00;
            14'd7202: data <= 8'h00;
            14'd7203: data <= 8'h00;
            14'd7204: data <= 8'h00;
            14'd7205: data <= 8'h00;
            14'd7206: data <= 8'h0F;
            14'd7207: data <= 8'hFF;
            14'd7208: data <= 8'hFF;
            14'd7209: data <= 8'hFF;
            14'd7210: data <= 8'hFF;
            14'd7211: data <= 8'hFF;
            14'd7212: data <= 8'hFF;
            14'd7213: data <= 8'hFF;
            14'd7214: data <= 8'hFF;
            14'd7215: data <= 8'hFF;
            14'd7216: data <= 8'hFF;
            14'd7217: data <= 8'hFF;
            14'd7218: data <= 8'hFF;
            14'd7219: data <= 8'hFF;
            14'd7220: data <= 8'hFF;
            14'd7221: data <= 8'hFF;
            14'd7222: data <= 8'hFF;
            14'd7223: data <= 8'hFF;
            14'd7224: data <= 8'hFF;
            14'd7225: data <= 8'hFF;
            14'd7226: data <= 8'hFF;
            14'd7227: data <= 8'hFF;
            14'd7228: data <= 8'hFF;
            14'd7229: data <= 8'hFF;
            14'd7230: data <= 8'hFF;
            14'd7231: data <= 8'hFF;
            14'd7232: data <= 8'hFF;
            14'd7233: data <= 8'hF0;
            14'd7234: data <= 8'h00;
            14'd7235: data <= 8'h00;
            14'd7236: data <= 8'h00;
            14'd7237: data <= 8'h00;
            14'd7238: data <= 8'h00;
            14'd7239: data <= 8'h00;
            14'd7240: data <= 8'h00;
            14'd7241: data <= 8'h00;
            14'd7242: data <= 8'h00;
            14'd7243: data <= 8'h00;
            14'd7244: data <= 8'h00;
            14'd7245: data <= 8'h00;
            14'd7246: data <= 8'h0F;
            14'd7247: data <= 8'hFF;
            14'd7248: data <= 8'hFF;
            14'd7249: data <= 8'hFF;
            14'd7250: data <= 8'hFF;
            14'd7251: data <= 8'hFF;
            14'd7252: data <= 8'hFF;
            14'd7253: data <= 8'hFF;
            14'd7254: data <= 8'hFF;
            14'd7255: data <= 8'hFF;
            14'd7256: data <= 8'hFF;
            14'd7257: data <= 8'hFF;
            14'd7258: data <= 8'hFF;
            14'd7259: data <= 8'hFF;
            14'd7260: data <= 8'hFF;
            14'd7261: data <= 8'hFF;
            14'd7262: data <= 8'hFF;
            14'd7263: data <= 8'hFF;
            14'd7264: data <= 8'hFF;
            14'd7265: data <= 8'hFF;
            14'd7266: data <= 8'hFF;
            14'd7267: data <= 8'hFF;
            14'd7268: data <= 8'hFF;
            14'd7269: data <= 8'hFF;
            14'd7270: data <= 8'hFF;
            14'd7271: data <= 8'hFF;
            14'd7272: data <= 8'hFF;
            14'd7273: data <= 8'hF0;
            14'd7274: data <= 8'h00;
            14'd7275: data <= 8'h00;
            14'd7276: data <= 8'h00;
            14'd7277: data <= 8'h00;
            14'd7278: data <= 8'h00;
            14'd7279: data <= 8'h00;
            14'd7280: data <= 8'h00;
            14'd7281: data <= 8'h00;
            14'd7282: data <= 8'h00;
            14'd7283: data <= 8'h00;
            14'd7284: data <= 8'h00;
            14'd7285: data <= 8'h00;
            14'd7286: data <= 8'h0F;
            14'd7287: data <= 8'hFF;
            14'd7288: data <= 8'hFF;
            14'd7289: data <= 8'hFF;
            14'd7290: data <= 8'hFF;
            14'd7291: data <= 8'hFF;
            14'd7292: data <= 8'hFF;
            14'd7293: data <= 8'hFF;
            14'd7294: data <= 8'hFF;
            14'd7295: data <= 8'hFF;
            14'd7296: data <= 8'hFF;
            14'd7297: data <= 8'hFF;
            14'd7298: data <= 8'hFF;
            14'd7299: data <= 8'hFF;
            14'd7300: data <= 8'hFF;
            14'd7301: data <= 8'hFF;
            14'd7302: data <= 8'hFF;
            14'd7303: data <= 8'hFF;
            14'd7304: data <= 8'hFF;
            14'd7305: data <= 8'hFF;
            14'd7306: data <= 8'hFF;
            14'd7307: data <= 8'hFF;
            14'd7308: data <= 8'hFF;
            14'd7309: data <= 8'hFF;
            14'd7310: data <= 8'hFF;
            14'd7311: data <= 8'hFF;
            14'd7312: data <= 8'hFF;
            14'd7313: data <= 8'hF0;
            14'd7314: data <= 8'h00;
            14'd7315: data <= 8'h00;
            14'd7316: data <= 8'h00;
            14'd7317: data <= 8'h00;
            14'd7318: data <= 8'h00;
            14'd7319: data <= 8'h00;
            14'd7320: data <= 8'h00;
            14'd7321: data <= 8'h00;
            14'd7322: data <= 8'h00;
            14'd7323: data <= 8'h00;
            14'd7324: data <= 8'h00;
            14'd7325: data <= 8'h00;
            14'd7326: data <= 8'h0F;
            14'd7327: data <= 8'hFF;
            14'd7328: data <= 8'hFF;
            14'd7329: data <= 8'hFF;
            14'd7330: data <= 8'hFF;
            14'd7331: data <= 8'hFF;
            14'd7332: data <= 8'hFF;
            14'd7333: data <= 8'hFF;
            14'd7334: data <= 8'hBF;
            14'd7335: data <= 8'hFF;
            14'd7336: data <= 8'hFF;
            14'd7337: data <= 8'hFF;
            14'd7338: data <= 8'hFF;
            14'd7339: data <= 8'hFF;
            14'd7340: data <= 8'hFF;
            14'd7341: data <= 8'hFF;
            14'd7342: data <= 8'hFF;
            14'd7343: data <= 8'hFF;
            14'd7344: data <= 8'hFF;
            14'd7345: data <= 8'hFF;
            14'd7346: data <= 8'hFF;
            14'd7347: data <= 8'hFF;
            14'd7348: data <= 8'hFF;
            14'd7349: data <= 8'hFF;
            14'd7350: data <= 8'hFF;
            14'd7351: data <= 8'hFF;
            14'd7352: data <= 8'hFF;
            14'd7353: data <= 8'hF0;
            14'd7354: data <= 8'h00;
            14'd7355: data <= 8'h00;
            14'd7356: data <= 8'h00;
            14'd7357: data <= 8'h00;
            14'd7358: data <= 8'h00;
            14'd7359: data <= 8'h00;
            14'd7360: data <= 8'h00;
            14'd7361: data <= 8'h00;
            14'd7362: data <= 8'h00;
            14'd7363: data <= 8'h00;
            14'd7364: data <= 8'h00;
            14'd7365: data <= 8'h00;
            14'd7366: data <= 8'h0F;
            14'd7367: data <= 8'hFF;
            14'd7368: data <= 8'hFF;
            14'd7369: data <= 8'hFF;
            14'd7370: data <= 8'hFF;
            14'd7371: data <= 8'hFF;
            14'd7372: data <= 8'hFF;
            14'd7373: data <= 8'hFF;
            14'd7374: data <= 8'hFF;
            14'd7375: data <= 8'hFF;
            14'd7376: data <= 8'hFF;
            14'd7377: data <= 8'hFF;
            14'd7378: data <= 8'hFF;
            14'd7379: data <= 8'hFF;
            14'd7380: data <= 8'hFF;
            14'd7381: data <= 8'hFF;
            14'd7382: data <= 8'hFF;
            14'd7383: data <= 8'hFF;
            14'd7384: data <= 8'hFF;
            14'd7385: data <= 8'hFF;
            14'd7386: data <= 8'hFF;
            14'd7387: data <= 8'hFF;
            14'd7388: data <= 8'hFF;
            14'd7389: data <= 8'hFF;
            14'd7390: data <= 8'hFF;
            14'd7391: data <= 8'hFF;
            14'd7392: data <= 8'hFF;
            14'd7393: data <= 8'hF0;
            14'd7394: data <= 8'h00;
            14'd7395: data <= 8'h00;
            14'd7396: data <= 8'h00;
            14'd7397: data <= 8'h00;
            14'd7398: data <= 8'h00;
            14'd7399: data <= 8'h00;
            14'd7400: data <= 8'h00;
            14'd7401: data <= 8'h00;
            14'd7402: data <= 8'h00;
            14'd7403: data <= 8'h00;
            14'd7404: data <= 8'h00;
            14'd7405: data <= 8'h00;
            14'd7406: data <= 8'h0F;
            14'd7407: data <= 8'hFF;
            14'd7408: data <= 8'hFF;
            14'd7409: data <= 8'hFF;
            14'd7410: data <= 8'hFF;
            14'd7411: data <= 8'hFF;
            14'd7412: data <= 8'hFF;
            14'd7413: data <= 8'hFF;
            14'd7414: data <= 8'hFF;
            14'd7415: data <= 8'hFF;
            14'd7416: data <= 8'hFF;
            14'd7417: data <= 8'hFF;
            14'd7418: data <= 8'hFF;
            14'd7419: data <= 8'hFF;
            14'd7420: data <= 8'hFF;
            14'd7421: data <= 8'hFE;
            14'd7422: data <= 8'hFF;
            14'd7423: data <= 8'hFF;
            14'd7424: data <= 8'hFF;
            14'd7425: data <= 8'hFF;
            14'd7426: data <= 8'hFF;
            14'd7427: data <= 8'hFF;
            14'd7428: data <= 8'hFF;
            14'd7429: data <= 8'hFF;
            14'd7430: data <= 8'hFF;
            14'd7431: data <= 8'hFF;
            14'd7432: data <= 8'hFF;
            14'd7433: data <= 8'hF0;
            14'd7434: data <= 8'h00;
            14'd7435: data <= 8'h00;
            14'd7436: data <= 8'h00;
            14'd7437: data <= 8'h00;
            14'd7438: data <= 8'h00;
            14'd7439: data <= 8'h00;
            14'd7440: data <= 8'h00;
            14'd7441: data <= 8'h00;
            14'd7442: data <= 8'h00;
            14'd7443: data <= 8'h00;
            14'd7444: data <= 8'h00;
            14'd7445: data <= 8'h00;
            14'd7446: data <= 8'h0F;
            14'd7447: data <= 8'hFF;
            14'd7448: data <= 8'hFF;
            14'd7449: data <= 8'hFF;
            14'd7450: data <= 8'hFF;
            14'd7451: data <= 8'hFF;
            14'd7452: data <= 8'hFF;
            14'd7453: data <= 8'hFF;
            14'd7454: data <= 8'hFF;
            14'd7455: data <= 8'hFF;
            14'd7456: data <= 8'hFF;
            14'd7457: data <= 8'hFF;
            14'd7458: data <= 8'hFF;
            14'd7459: data <= 8'hFF;
            14'd7460: data <= 8'hFF;
            14'd7461: data <= 8'hFF;
            14'd7462: data <= 8'hFF;
            14'd7463: data <= 8'hFF;
            14'd7464: data <= 8'hFF;
            14'd7465: data <= 8'hFF;
            14'd7466: data <= 8'hFF;
            14'd7467: data <= 8'hFF;
            14'd7468: data <= 8'hFF;
            14'd7469: data <= 8'hFF;
            14'd7470: data <= 8'hFF;
            14'd7471: data <= 8'hFF;
            14'd7472: data <= 8'hFF;
            14'd7473: data <= 8'hF0;
            14'd7474: data <= 8'h00;
            14'd7475: data <= 8'h00;
            14'd7476: data <= 8'h00;
            14'd7477: data <= 8'h00;
            14'd7478: data <= 8'h00;
            14'd7479: data <= 8'h00;
            14'd7480: data <= 8'h00;
            14'd7481: data <= 8'h00;
            14'd7482: data <= 8'h00;
            14'd7483: data <= 8'h00;
            14'd7484: data <= 8'h00;
            14'd7485: data <= 8'h00;
            14'd7486: data <= 8'h0F;
            14'd7487: data <= 8'hFF;
            14'd7488: data <= 8'hFF;
            14'd7489: data <= 8'hFF;
            14'd7490: data <= 8'hFF;
            14'd7491: data <= 8'hFF;
            14'd7492: data <= 8'hFF;
            14'd7493: data <= 8'hFF;
            14'd7494: data <= 8'hFF;
            14'd7495: data <= 8'hFF;
            14'd7496: data <= 8'hFF;
            14'd7497: data <= 8'hFF;
            14'd7498: data <= 8'hFF;
            14'd7499: data <= 8'hFF;
            14'd7500: data <= 8'hFF;
            14'd7501: data <= 8'hFF;
            14'd7502: data <= 8'hFF;
            14'd7503: data <= 8'hFF;
            14'd7504: data <= 8'hFF;
            14'd7505: data <= 8'hFF;
            14'd7506: data <= 8'hFF;
            14'd7507: data <= 8'hFF;
            14'd7508: data <= 8'hFF;
            14'd7509: data <= 8'hFF;
            14'd7510: data <= 8'hFF;
            14'd7511: data <= 8'hFF;
            14'd7512: data <= 8'hFF;
            14'd7513: data <= 8'hF0;
            14'd7514: data <= 8'h00;
            14'd7515: data <= 8'h00;
            14'd7516: data <= 8'h00;
            14'd7517: data <= 8'h00;
            14'd7518: data <= 8'h00;
            14'd7519: data <= 8'h00;
            14'd7520: data <= 8'h00;
            14'd7521: data <= 8'h00;
            14'd7522: data <= 8'h00;
            14'd7523: data <= 8'h00;
            14'd7524: data <= 8'h00;
            14'd7525: data <= 8'h00;
            14'd7526: data <= 8'h0F;
            14'd7527: data <= 8'hFF;
            14'd7528: data <= 8'hFF;
            14'd7529: data <= 8'hFF;
            14'd7530: data <= 8'hFF;
            14'd7531: data <= 8'hFF;
            14'd7532: data <= 8'hFF;
            14'd7533: data <= 8'hFF;
            14'd7534: data <= 8'hFF;
            14'd7535: data <= 8'hFF;
            14'd7536: data <= 8'hFF;
            14'd7537: data <= 8'hFF;
            14'd7538: data <= 8'hFF;
            14'd7539: data <= 8'hFF;
            14'd7540: data <= 8'hFF;
            14'd7541: data <= 8'hFF;
            14'd7542: data <= 8'hFF;
            14'd7543: data <= 8'hFF;
            14'd7544: data <= 8'hFF;
            14'd7545: data <= 8'hFF;
            14'd7546: data <= 8'hFF;
            14'd7547: data <= 8'hFF;
            14'd7548: data <= 8'hFF;
            14'd7549: data <= 8'hFF;
            14'd7550: data <= 8'hFF;
            14'd7551: data <= 8'hFF;
            14'd7552: data <= 8'hFF;
            14'd7553: data <= 8'hF0;
            14'd7554: data <= 8'h00;
            14'd7555: data <= 8'h00;
            14'd7556: data <= 8'h00;
            14'd7557: data <= 8'h00;
            14'd7558: data <= 8'h00;
            14'd7559: data <= 8'h00;
            14'd7560: data <= 8'h00;
            14'd7561: data <= 8'h00;
            14'd7562: data <= 8'h00;
            14'd7563: data <= 8'h00;
            14'd7564: data <= 8'h00;
            14'd7565: data <= 8'h00;
            14'd7566: data <= 8'h0F;
            14'd7567: data <= 8'hFF;
            14'd7568: data <= 8'hFF;
            14'd7569: data <= 8'hFF;
            14'd7570: data <= 8'hFF;
            14'd7571: data <= 8'hFF;
            14'd7572: data <= 8'hFF;
            14'd7573: data <= 8'hFF;
            14'd7574: data <= 8'hFF;
            14'd7575: data <= 8'hFF;
            14'd7576: data <= 8'hFF;
            14'd7577: data <= 8'hFF;
            14'd7578: data <= 8'hFF;
            14'd7579: data <= 8'hFF;
            14'd7580: data <= 8'hFF;
            14'd7581: data <= 8'hFF;
            14'd7582: data <= 8'hFF;
            14'd7583: data <= 8'hFF;
            14'd7584: data <= 8'hFF;
            14'd7585: data <= 8'hFF;
            14'd7586: data <= 8'hFF;
            14'd7587: data <= 8'hFF;
            14'd7588: data <= 8'hFF;
            14'd7589: data <= 8'hFF;
            14'd7590: data <= 8'hFF;
            14'd7591: data <= 8'hFF;
            14'd7592: data <= 8'hFF;
            14'd7593: data <= 8'hF0;
            14'd7594: data <= 8'h00;
            14'd7595: data <= 8'h00;
            14'd7596: data <= 8'h00;
            14'd7597: data <= 8'h00;
            14'd7598: data <= 8'h00;
            14'd7599: data <= 8'h00;
            14'd7600: data <= 8'h00;
            14'd7601: data <= 8'h00;
            14'd7602: data <= 8'h00;
            14'd7603: data <= 8'h00;
            14'd7604: data <= 8'h00;
            14'd7605: data <= 8'h00;
            14'd7606: data <= 8'h0F;
            14'd7607: data <= 8'hFF;
            14'd7608: data <= 8'hFF;
            14'd7609: data <= 8'hFF;
            14'd7610: data <= 8'hFF;
            14'd7611: data <= 8'hFF;
            14'd7612: data <= 8'hFF;
            14'd7613: data <= 8'hFF;
            14'd7614: data <= 8'hFF;
            14'd7615: data <= 8'hFF;
            14'd7616: data <= 8'hFF;
            14'd7617: data <= 8'hFF;
            14'd7618: data <= 8'hFF;
            14'd7619: data <= 8'hFF;
            14'd7620: data <= 8'hFF;
            14'd7621: data <= 8'hFF;
            14'd7622: data <= 8'hFF;
            14'd7623: data <= 8'hFF;
            14'd7624: data <= 8'hFF;
            14'd7625: data <= 8'hFF;
            14'd7626: data <= 8'hFF;
            14'd7627: data <= 8'hFF;
            14'd7628: data <= 8'hFF;
            14'd7629: data <= 8'hFF;
            14'd7630: data <= 8'hFF;
            14'd7631: data <= 8'hFF;
            14'd7632: data <= 8'hFF;
            14'd7633: data <= 8'hF0;
            14'd7634: data <= 8'h00;
            14'd7635: data <= 8'h00;
            14'd7636: data <= 8'h00;
            14'd7637: data <= 8'h00;
            14'd7638: data <= 8'h00;
            14'd7639: data <= 8'h00;
            14'd7640: data <= 8'h00;
            14'd7641: data <= 8'h00;
            14'd7642: data <= 8'h00;
            14'd7643: data <= 8'h00;
            14'd7644: data <= 8'h00;
            14'd7645: data <= 8'h00;
            14'd7646: data <= 8'h0F;
            14'd7647: data <= 8'hFF;
            14'd7648: data <= 8'hFF;
            14'd7649: data <= 8'hFF;
            14'd7650: data <= 8'hFF;
            14'd7651: data <= 8'hFF;
            14'd7652: data <= 8'hFF;
            14'd7653: data <= 8'hFF;
            14'd7654: data <= 8'hFF;
            14'd7655: data <= 8'hFF;
            14'd7656: data <= 8'hFF;
            14'd7657: data <= 8'hFF;
            14'd7658: data <= 8'hFF;
            14'd7659: data <= 8'hFF;
            14'd7660: data <= 8'hFF;
            14'd7661: data <= 8'hFF;
            14'd7662: data <= 8'hFF;
            14'd7663: data <= 8'hFF;
            14'd7664: data <= 8'hFF;
            14'd7665: data <= 8'hFF;
            14'd7666: data <= 8'hFF;
            14'd7667: data <= 8'hFF;
            14'd7668: data <= 8'hFF;
            14'd7669: data <= 8'hFF;
            14'd7670: data <= 8'hFF;
            14'd7671: data <= 8'hFF;
            14'd7672: data <= 8'hFF;
            14'd7673: data <= 8'hF0;
            14'd7674: data <= 8'h00;
            14'd7675: data <= 8'h00;
            14'd7676: data <= 8'h00;
            14'd7677: data <= 8'h00;
            14'd7678: data <= 8'h00;
            14'd7679: data <= 8'h00;
            14'd7680: data <= 8'h00;
            14'd7681: data <= 8'h00;
            14'd7682: data <= 8'h00;
            14'd7683: data <= 8'h00;
            14'd7684: data <= 8'h00;
            14'd7685: data <= 8'h00;
            14'd7686: data <= 8'h0F;
            14'd7687: data <= 8'hFF;
            14'd7688: data <= 8'hFF;
            14'd7689: data <= 8'hFF;
            14'd7690: data <= 8'hFF;
            14'd7691: data <= 8'hFF;
            14'd7692: data <= 8'hFF;
            14'd7693: data <= 8'hFF;
            14'd7694: data <= 8'hFF;
            14'd7695: data <= 8'hFF;
            14'd7696: data <= 8'hFF;
            14'd7697: data <= 8'hFE;
            14'd7698: data <= 8'hFF;
            14'd7699: data <= 8'hFF;
            14'd7700: data <= 8'hF8;
            14'd7701: data <= 8'hFF;
            14'd7702: data <= 8'hFF;
            14'd7703: data <= 8'hFF;
            14'd7704: data <= 8'hFF;
            14'd7705: data <= 8'hFF;
            14'd7706: data <= 8'hFF;
            14'd7707: data <= 8'hFF;
            14'd7708: data <= 8'hFF;
            14'd7709: data <= 8'hFF;
            14'd7710: data <= 8'hFF;
            14'd7711: data <= 8'hFF;
            14'd7712: data <= 8'hFF;
            14'd7713: data <= 8'hF0;
            14'd7714: data <= 8'h00;
            14'd7715: data <= 8'h00;
            14'd7716: data <= 8'h00;
            14'd7717: data <= 8'h00;
            14'd7718: data <= 8'h00;
            14'd7719: data <= 8'h00;
            14'd7720: data <= 8'h00;
            14'd7721: data <= 8'h00;
            14'd7722: data <= 8'h00;
            14'd7723: data <= 8'h00;
            14'd7724: data <= 8'h00;
            14'd7725: data <= 8'h00;
            14'd7726: data <= 8'h0F;
            14'd7727: data <= 8'hFF;
            14'd7728: data <= 8'hFF;
            14'd7729: data <= 8'hFF;
            14'd7730: data <= 8'hFF;
            14'd7731: data <= 8'hFF;
            14'd7732: data <= 8'hFF;
            14'd7733: data <= 8'hFF;
            14'd7734: data <= 8'hFF;
            14'd7735: data <= 8'hFF;
            14'd7736: data <= 8'hFF;
            14'd7737: data <= 8'hBC;
            14'd7738: data <= 8'h7F;
            14'd7739: data <= 8'hFF;
            14'd7740: data <= 8'hF8;
            14'd7741: data <= 8'h72;
            14'd7742: data <= 8'h7F;
            14'd7743: data <= 8'hFF;
            14'd7744: data <= 8'hFF;
            14'd7745: data <= 8'hFF;
            14'd7746: data <= 8'hFF;
            14'd7747: data <= 8'hFF;
            14'd7748: data <= 8'hFF;
            14'd7749: data <= 8'hFF;
            14'd7750: data <= 8'hFF;
            14'd7751: data <= 8'hFF;
            14'd7752: data <= 8'hFF;
            14'd7753: data <= 8'hF0;
            14'd7754: data <= 8'h00;
            14'd7755: data <= 8'h00;
            14'd7756: data <= 8'h00;
            14'd7757: data <= 8'h00;
            14'd7758: data <= 8'h00;
            14'd7759: data <= 8'h00;
            14'd7760: data <= 8'h00;
            14'd7761: data <= 8'h00;
            14'd7762: data <= 8'h00;
            14'd7763: data <= 8'h00;
            14'd7764: data <= 8'h00;
            14'd7765: data <= 8'h00;
            14'd7766: data <= 8'h0F;
            14'd7767: data <= 8'hFF;
            14'd7768: data <= 8'hFF;
            14'd7769: data <= 8'hFF;
            14'd7770: data <= 8'hFF;
            14'd7771: data <= 8'hFF;
            14'd7772: data <= 8'hFF;
            14'd7773: data <= 8'hFF;
            14'd7774: data <= 8'hFF;
            14'd7775: data <= 8'hFF;
            14'd7776: data <= 8'hFF;
            14'd7777: data <= 8'h18;
            14'd7778: data <= 8'h7F;
            14'd7779: data <= 8'hFF;
            14'd7780: data <= 8'hF8;
            14'd7781: data <= 8'h00;
            14'd7782: data <= 8'h1F;
            14'd7783: data <= 8'hFF;
            14'd7784: data <= 8'hFF;
            14'd7785: data <= 8'hFF;
            14'd7786: data <= 8'hFF;
            14'd7787: data <= 8'hFF;
            14'd7788: data <= 8'hFF;
            14'd7789: data <= 8'hFF;
            14'd7790: data <= 8'hFF;
            14'd7791: data <= 8'hFF;
            14'd7792: data <= 8'hFF;
            14'd7793: data <= 8'hF0;
            14'd7794: data <= 8'h00;
            14'd7795: data <= 8'h00;
            14'd7796: data <= 8'h00;
            14'd7797: data <= 8'h00;
            14'd7798: data <= 8'h00;
            14'd7799: data <= 8'h00;
            14'd7800: data <= 8'h00;
            14'd7801: data <= 8'h00;
            14'd7802: data <= 8'h00;
            14'd7803: data <= 8'h00;
            14'd7804: data <= 8'h00;
            14'd7805: data <= 8'h00;
            14'd7806: data <= 8'h0F;
            14'd7807: data <= 8'hFF;
            14'd7808: data <= 8'hFF;
            14'd7809: data <= 8'hFF;
            14'd7810: data <= 8'hFF;
            14'd7811: data <= 8'hFF;
            14'd7812: data <= 8'hFF;
            14'd7813: data <= 8'hFF;
            14'd7814: data <= 8'hFF;
            14'd7815: data <= 8'hFF;
            14'd7816: data <= 8'hFF;
            14'd7817: data <= 8'h08;
            14'd7818: data <= 8'h7F;
            14'd7819: data <= 8'hFF;
            14'd7820: data <= 8'hF0;
            14'd7821: data <= 8'h00;
            14'd7822: data <= 8'h0F;
            14'd7823: data <= 8'hFF;
            14'd7824: data <= 8'hFF;
            14'd7825: data <= 8'hFF;
            14'd7826: data <= 8'hFF;
            14'd7827: data <= 8'hFF;
            14'd7828: data <= 8'hFF;
            14'd7829: data <= 8'hFF;
            14'd7830: data <= 8'hFF;
            14'd7831: data <= 8'hFF;
            14'd7832: data <= 8'hFF;
            14'd7833: data <= 8'hF0;
            14'd7834: data <= 8'h00;
            14'd7835: data <= 8'h00;
            14'd7836: data <= 8'h00;
            14'd7837: data <= 8'h00;
            14'd7838: data <= 8'h00;
            14'd7839: data <= 8'h00;
            14'd7840: data <= 8'h00;
            14'd7841: data <= 8'h00;
            14'd7842: data <= 8'h00;
            14'd7843: data <= 8'h00;
            14'd7844: data <= 8'h00;
            14'd7845: data <= 8'h00;
            14'd7846: data <= 8'h0F;
            14'd7847: data <= 8'hFF;
            14'd7848: data <= 8'hFF;
            14'd7849: data <= 8'hFF;
            14'd7850: data <= 8'hFF;
            14'd7851: data <= 8'hFF;
            14'd7852: data <= 8'hFF;
            14'd7853: data <= 8'hFF;
            14'd7854: data <= 8'hFF;
            14'd7855: data <= 8'hFF;
            14'd7856: data <= 8'hFF;
            14'd7857: data <= 8'h18;
            14'd7858: data <= 8'h03;
            14'd7859: data <= 8'hFF;
            14'd7860: data <= 8'hF0;
            14'd7861: data <= 8'h00;
            14'd7862: data <= 8'h1F;
            14'd7863: data <= 8'hFF;
            14'd7864: data <= 8'hF8;
            14'd7865: data <= 8'h7F;
            14'd7866: data <= 8'hFF;
            14'd7867: data <= 8'hFF;
            14'd7868: data <= 8'hFF;
            14'd7869: data <= 8'hFF;
            14'd7870: data <= 8'hFF;
            14'd7871: data <= 8'hFF;
            14'd7872: data <= 8'hFF;
            14'd7873: data <= 8'hF0;
            14'd7874: data <= 8'h00;
            14'd7875: data <= 8'h00;
            14'd7876: data <= 8'h00;
            14'd7877: data <= 8'h00;
            14'd7878: data <= 8'h00;
            14'd7879: data <= 8'h00;
            14'd7880: data <= 8'h00;
            14'd7881: data <= 8'h00;
            14'd7882: data <= 8'h00;
            14'd7883: data <= 8'h00;
            14'd7884: data <= 8'h00;
            14'd7885: data <= 8'h00;
            14'd7886: data <= 8'h0F;
            14'd7887: data <= 8'hFF;
            14'd7888: data <= 8'hFF;
            14'd7889: data <= 8'hFF;
            14'd7890: data <= 8'hFF;
            14'd7891: data <= 8'hFF;
            14'd7892: data <= 8'hFF;
            14'd7893: data <= 8'hFF;
            14'd7894: data <= 8'hFF;
            14'd7895: data <= 8'hFF;
            14'd7896: data <= 8'hFE;
            14'd7897: data <= 8'h00;
            14'd7898: data <= 8'h01;
            14'd7899: data <= 8'hFF;
            14'd7900: data <= 8'hE1;
            14'd7901: data <= 8'hFF;
            14'd7902: data <= 8'hFF;
            14'd7903: data <= 8'hFF;
            14'd7904: data <= 8'hF8;
            14'd7905: data <= 8'h7F;
            14'd7906: data <= 8'hFF;
            14'd7907: data <= 8'hFF;
            14'd7908: data <= 8'hFF;
            14'd7909: data <= 8'hFF;
            14'd7910: data <= 8'hFF;
            14'd7911: data <= 8'hFF;
            14'd7912: data <= 8'hFF;
            14'd7913: data <= 8'hF0;
            14'd7914: data <= 8'h00;
            14'd7915: data <= 8'h00;
            14'd7916: data <= 8'h00;
            14'd7917: data <= 8'h00;
            14'd7918: data <= 8'h00;
            14'd7919: data <= 8'h00;
            14'd7920: data <= 8'h00;
            14'd7921: data <= 8'h00;
            14'd7922: data <= 8'h00;
            14'd7923: data <= 8'h00;
            14'd7924: data <= 8'h00;
            14'd7925: data <= 8'h00;
            14'd7926: data <= 8'h0F;
            14'd7927: data <= 8'hFF;
            14'd7928: data <= 8'hFF;
            14'd7929: data <= 8'hFF;
            14'd7930: data <= 8'hFF;
            14'd7931: data <= 8'hFF;
            14'd7932: data <= 8'hFF;
            14'd7933: data <= 8'hFF;
            14'd7934: data <= 8'hFF;
            14'd7935: data <= 8'hFF;
            14'd7936: data <= 8'hFE;
            14'd7937: data <= 8'h00;
            14'd7938: data <= 8'h03;
            14'd7939: data <= 8'hFF;
            14'd7940: data <= 8'hE3;
            14'd7941: data <= 8'hFE;
            14'd7942: data <= 8'h3F;
            14'd7943: data <= 8'hFF;
            14'd7944: data <= 8'hF8;
            14'd7945: data <= 8'h7F;
            14'd7946: data <= 8'hFF;
            14'd7947: data <= 8'hF7;
            14'd7948: data <= 8'hFF;
            14'd7949: data <= 8'hFF;
            14'd7950: data <= 8'hFF;
            14'd7951: data <= 8'hFF;
            14'd7952: data <= 8'hFF;
            14'd7953: data <= 8'hF0;
            14'd7954: data <= 8'h00;
            14'd7955: data <= 8'h00;
            14'd7956: data <= 8'h00;
            14'd7957: data <= 8'h00;
            14'd7958: data <= 8'h00;
            14'd7959: data <= 8'h00;
            14'd7960: data <= 8'h00;
            14'd7961: data <= 8'h00;
            14'd7962: data <= 8'h00;
            14'd7963: data <= 8'h00;
            14'd7964: data <= 8'h00;
            14'd7965: data <= 8'h00;
            14'd7966: data <= 8'h0F;
            14'd7967: data <= 8'hFF;
            14'd7968: data <= 8'hFF;
            14'd7969: data <= 8'hFF;
            14'd7970: data <= 8'hFF;
            14'd7971: data <= 8'hFF;
            14'd7972: data <= 8'hFF;
            14'd7973: data <= 8'hFF;
            14'd7974: data <= 8'hFF;
            14'd7975: data <= 8'hFF;
            14'd7976: data <= 8'hFE;
            14'd7977: data <= 8'h00;
            14'd7978: data <= 8'h03;
            14'd7979: data <= 8'hFF;
            14'd7980: data <= 8'hC4;
            14'd7981: data <= 8'h00;
            14'd7982: data <= 8'h1F;
            14'd7983: data <= 8'hFF;
            14'd7984: data <= 8'hF0;
            14'd7985: data <= 8'h7F;
            14'd7986: data <= 8'hFF;
            14'd7987: data <= 8'hFF;
            14'd7988: data <= 8'hFF;
            14'd7989: data <= 8'hFF;
            14'd7990: data <= 8'hFF;
            14'd7991: data <= 8'hFF;
            14'd7992: data <= 8'hFF;
            14'd7993: data <= 8'hF0;
            14'd7994: data <= 8'h00;
            14'd7995: data <= 8'h00;
            14'd7996: data <= 8'h00;
            14'd7997: data <= 8'h00;
            14'd7998: data <= 8'h00;
            14'd7999: data <= 8'h00;
            14'd8000: data <= 8'h00;
            14'd8001: data <= 8'h00;
            14'd8002: data <= 8'h00;
            14'd8003: data <= 8'h00;
            14'd8004: data <= 8'h00;
            14'd8005: data <= 8'h00;
            14'd8006: data <= 8'h0F;
            14'd8007: data <= 8'hFF;
            14'd8008: data <= 8'hFF;
            14'd8009: data <= 8'hFF;
            14'd8010: data <= 8'hFF;
            14'd8011: data <= 8'hFF;
            14'd8012: data <= 8'hFF;
            14'd8013: data <= 8'hFF;
            14'd8014: data <= 8'hFF;
            14'd8015: data <= 8'hFF;
            14'd8016: data <= 8'hFC;
            14'd8017: data <= 8'h18;
            14'd8018: data <= 8'h7F;
            14'd8019: data <= 8'hFF;
            14'd8020: data <= 8'h84;
            14'd8021: data <= 8'h00;
            14'd8022: data <= 8'h3F;
            14'd8023: data <= 8'hFF;
            14'd8024: data <= 8'hF8;
            14'd8025: data <= 8'h7F;
            14'd8026: data <= 8'hFF;
            14'd8027: data <= 8'hFF;
            14'd8028: data <= 8'hFF;
            14'd8029: data <= 8'hFF;
            14'd8030: data <= 8'hFF;
            14'd8031: data <= 8'hFF;
            14'd8032: data <= 8'hFF;
            14'd8033: data <= 8'hF0;
            14'd8034: data <= 8'h00;
            14'd8035: data <= 8'h00;
            14'd8036: data <= 8'h00;
            14'd8037: data <= 8'h00;
            14'd8038: data <= 8'h00;
            14'd8039: data <= 8'h00;
            14'd8040: data <= 8'h00;
            14'd8041: data <= 8'h00;
            14'd8042: data <= 8'h00;
            14'd8043: data <= 8'h00;
            14'd8044: data <= 8'h00;
            14'd8045: data <= 8'h00;
            14'd8046: data <= 8'h0F;
            14'd8047: data <= 8'hFF;
            14'd8048: data <= 8'hFF;
            14'd8049: data <= 8'hFF;
            14'd8050: data <= 8'hFF;
            14'd8051: data <= 8'hFF;
            14'd8052: data <= 8'hFF;
            14'd8053: data <= 8'hFF;
            14'd8054: data <= 8'hFF;
            14'd8055: data <= 8'hFF;
            14'd8056: data <= 8'hF8;
            14'd8057: data <= 8'h38;
            14'd8058: data <= 8'h7F;
            14'd8059: data <= 8'hFF;
            14'd8060: data <= 8'h8C;
            14'd8061: data <= 8'h3E;
            14'd8062: data <= 8'h7F;
            14'd8063: data <= 8'hFF;
            14'd8064: data <= 8'hF0;
            14'd8065: data <= 8'hFF;
            14'd8066: data <= 8'hFF;
            14'd8067: data <= 8'hFF;
            14'd8068: data <= 8'hFF;
            14'd8069: data <= 8'hFF;
            14'd8070: data <= 8'hFF;
            14'd8071: data <= 8'hFF;
            14'd8072: data <= 8'hFF;
            14'd8073: data <= 8'hF0;
            14'd8074: data <= 8'h00;
            14'd8075: data <= 8'h00;
            14'd8076: data <= 8'h00;
            14'd8077: data <= 8'h00;
            14'd8078: data <= 8'h00;
            14'd8079: data <= 8'h00;
            14'd8080: data <= 8'h00;
            14'd8081: data <= 8'h00;
            14'd8082: data <= 8'h00;
            14'd8083: data <= 8'h00;
            14'd8084: data <= 8'h00;
            14'd8085: data <= 8'h00;
            14'd8086: data <= 8'h0F;
            14'd8087: data <= 8'hFF;
            14'd8088: data <= 8'hFF;
            14'd8089: data <= 8'hFF;
            14'd8090: data <= 8'hFF;
            14'd8091: data <= 8'hFF;
            14'd8092: data <= 8'hFF;
            14'd8093: data <= 8'hFF;
            14'd8094: data <= 8'hFF;
            14'd8095: data <= 8'hFF;
            14'd8096: data <= 8'hE8;
            14'd8097: data <= 8'h78;
            14'd8098: data <= 8'h7F;
            14'd8099: data <= 8'hFF;
            14'd8100: data <= 8'hFF;
            14'd8101: data <= 8'h82;
            14'd8102: data <= 8'hDF;
            14'd8103: data <= 8'hFF;
            14'd8104: data <= 8'hF0;
            14'd8105: data <= 8'hFF;
            14'd8106: data <= 8'hFF;
            14'd8107: data <= 8'hFF;
            14'd8108: data <= 8'hFF;
            14'd8109: data <= 8'hFF;
            14'd8110: data <= 8'hFF;
            14'd8111: data <= 8'hFF;
            14'd8112: data <= 8'hFF;
            14'd8113: data <= 8'hF0;
            14'd8114: data <= 8'h00;
            14'd8115: data <= 8'h00;
            14'd8116: data <= 8'h00;
            14'd8117: data <= 8'h00;
            14'd8118: data <= 8'h00;
            14'd8119: data <= 8'h00;
            14'd8120: data <= 8'h00;
            14'd8121: data <= 8'h00;
            14'd8122: data <= 8'h00;
            14'd8123: data <= 8'h00;
            14'd8124: data <= 8'h00;
            14'd8125: data <= 8'h00;
            14'd8126: data <= 8'h0F;
            14'd8127: data <= 8'hFF;
            14'd8128: data <= 8'hFF;
            14'd8129: data <= 8'hFF;
            14'd8130: data <= 8'hFF;
            14'd8131: data <= 8'hFF;
            14'd8132: data <= 8'hFF;
            14'd8133: data <= 8'hFF;
            14'd8134: data <= 8'hFF;
            14'd8135: data <= 8'hFF;
            14'd8136: data <= 8'hF8;
            14'd8137: data <= 8'h7C;
            14'd8138: data <= 8'h7F;
            14'd8139: data <= 8'hFF;
            14'd8140: data <= 8'hFC;
            14'd8141: data <= 8'h00;
            14'd8142: data <= 8'h0F;
            14'd8143: data <= 8'hFF;
            14'd8144: data <= 8'hF0;
            14'd8145: data <= 8'h7F;
            14'd8146: data <= 8'hFF;
            14'd8147: data <= 8'hFF;
            14'd8148: data <= 8'hFF;
            14'd8149: data <= 8'hFF;
            14'd8150: data <= 8'hFF;
            14'd8151: data <= 8'hFF;
            14'd8152: data <= 8'hFF;
            14'd8153: data <= 8'hF0;
            14'd8154: data <= 8'h00;
            14'd8155: data <= 8'h00;
            14'd8156: data <= 8'h00;
            14'd8157: data <= 8'h00;
            14'd8158: data <= 8'h00;
            14'd8159: data <= 8'h00;
            14'd8160: data <= 8'h00;
            14'd8161: data <= 8'h00;
            14'd8162: data <= 8'h00;
            14'd8163: data <= 8'h00;
            14'd8164: data <= 8'h00;
            14'd8165: data <= 8'h00;
            14'd8166: data <= 8'h0F;
            14'd8167: data <= 8'hFF;
            14'd8168: data <= 8'hFF;
            14'd8169: data <= 8'hFF;
            14'd8170: data <= 8'hFF;
            14'd8171: data <= 8'hFF;
            14'd8172: data <= 8'hFF;
            14'd8173: data <= 8'hFF;
            14'd8174: data <= 8'hFF;
            14'd8175: data <= 8'hFF;
            14'd8176: data <= 8'hF8;
            14'd8177: data <= 8'hF8;
            14'd8178: data <= 8'h2F;
            14'd8179: data <= 8'hFF;
            14'd8180: data <= 8'hD8;
            14'd8181: data <= 8'h00;
            14'd8182: data <= 8'h0F;
            14'd8183: data <= 8'hFF;
            14'd8184: data <= 8'hF8;
            14'd8185: data <= 8'h7F;
            14'd8186: data <= 8'hFF;
            14'd8187: data <= 8'hFF;
            14'd8188: data <= 8'hFF;
            14'd8189: data <= 8'hFF;
            14'd8190: data <= 8'hFF;
            14'd8191: data <= 8'hFF;
            14'd8192: data <= 8'hFF;
            14'd8193: data <= 8'hF0;
            14'd8194: data <= 8'h00;
            14'd8195: data <= 8'h00;
            14'd8196: data <= 8'h00;
            14'd8197: data <= 8'h00;
            14'd8198: data <= 8'h00;
            14'd8199: data <= 8'h00;
            14'd8200: data <= 8'h00;
            14'd8201: data <= 8'h00;
            14'd8202: data <= 8'h00;
            14'd8203: data <= 8'h00;
            14'd8204: data <= 8'h00;
            14'd8205: data <= 8'h00;
            14'd8206: data <= 8'h0F;
            14'd8207: data <= 8'hFF;
            14'd8208: data <= 8'hFF;
            14'd8209: data <= 8'hFF;
            14'd8210: data <= 8'hFF;
            14'd8211: data <= 8'hFF;
            14'd8212: data <= 8'hFF;
            14'd8213: data <= 8'hFF;
            14'd8214: data <= 8'hFF;
            14'd8215: data <= 8'hFF;
            14'd8216: data <= 8'hFF;
            14'd8217: data <= 8'h80;
            14'd8218: data <= 8'h03;
            14'd8219: data <= 8'hFF;
            14'd8220: data <= 8'hFC;
            14'd8221: data <= 8'h00;
            14'd8222: data <= 8'h0F;
            14'd8223: data <= 8'hFF;
            14'd8224: data <= 8'hF8;
            14'd8225: data <= 8'hFF;
            14'd8226: data <= 8'hFF;
            14'd8227: data <= 8'hFF;
            14'd8228: data <= 8'hF7;
            14'd8229: data <= 8'hFF;
            14'd8230: data <= 8'hFF;
            14'd8231: data <= 8'hFF;
            14'd8232: data <= 8'hFF;
            14'd8233: data <= 8'hF0;
            14'd8234: data <= 8'h00;
            14'd8235: data <= 8'h00;
            14'd8236: data <= 8'h00;
            14'd8237: data <= 8'h00;
            14'd8238: data <= 8'h00;
            14'd8239: data <= 8'h00;
            14'd8240: data <= 8'h00;
            14'd8241: data <= 8'h00;
            14'd8242: data <= 8'h00;
            14'd8243: data <= 8'h00;
            14'd8244: data <= 8'h00;
            14'd8245: data <= 8'h00;
            14'd8246: data <= 8'h0F;
            14'd8247: data <= 8'hFF;
            14'd8248: data <= 8'hFF;
            14'd8249: data <= 8'hFF;
            14'd8250: data <= 8'hFF;
            14'd8251: data <= 8'hFF;
            14'd8252: data <= 8'hFF;
            14'd8253: data <= 8'hFF;
            14'd8254: data <= 8'hFF;
            14'd8255: data <= 8'hFF;
            14'd8256: data <= 8'hFF;
            14'd8257: data <= 8'h00;
            14'd8258: data <= 8'h03;
            14'd8259: data <= 8'hFF;
            14'd8260: data <= 8'hFF;
            14'd8261: data <= 8'hFF;
            14'd8262: data <= 8'h8F;
            14'd8263: data <= 8'hFF;
            14'd8264: data <= 8'hF8;
            14'd8265: data <= 8'hFF;
            14'd8266: data <= 8'hFF;
            14'd8267: data <= 8'hFF;
            14'd8268: data <= 8'hFF;
            14'd8269: data <= 8'hFF;
            14'd8270: data <= 8'hFF;
            14'd8271: data <= 8'hFF;
            14'd8272: data <= 8'hFF;
            14'd8273: data <= 8'hF0;
            14'd8274: data <= 8'h00;
            14'd8275: data <= 8'h00;
            14'd8276: data <= 8'h00;
            14'd8277: data <= 8'h00;
            14'd8278: data <= 8'h00;
            14'd8279: data <= 8'h00;
            14'd8280: data <= 8'h00;
            14'd8281: data <= 8'h00;
            14'd8282: data <= 8'h00;
            14'd8283: data <= 8'h00;
            14'd8284: data <= 8'h00;
            14'd8285: data <= 8'h00;
            14'd8286: data <= 8'h0F;
            14'd8287: data <= 8'hFF;
            14'd8288: data <= 8'hFF;
            14'd8289: data <= 8'hFF;
            14'd8290: data <= 8'hFF;
            14'd8291: data <= 8'hFF;
            14'd8292: data <= 8'hFF;
            14'd8293: data <= 8'hFF;
            14'd8294: data <= 8'hFF;
            14'd8295: data <= 8'hFF;
            14'd8296: data <= 8'hFF;
            14'd8297: data <= 8'h80;
            14'd8298: data <= 8'h03;
            14'd8299: data <= 8'hFF;
            14'd8300: data <= 8'hFF;
            14'd8301: data <= 8'hFF;
            14'd8302: data <= 8'h8F;
            14'd8303: data <= 8'hFF;
            14'd8304: data <= 8'hF9;
            14'd8305: data <= 8'hFF;
            14'd8306: data <= 8'hFF;
            14'd8307: data <= 8'hFF;
            14'd8308: data <= 8'hFF;
            14'd8309: data <= 8'hFF;
            14'd8310: data <= 8'hFF;
            14'd8311: data <= 8'hFF;
            14'd8312: data <= 8'hFF;
            14'd8313: data <= 8'hF0;
            14'd8314: data <= 8'h00;
            14'd8315: data <= 8'h00;
            14'd8316: data <= 8'h00;
            14'd8317: data <= 8'h00;
            14'd8318: data <= 8'h00;
            14'd8319: data <= 8'h00;
            14'd8320: data <= 8'h00;
            14'd8321: data <= 8'h00;
            14'd8322: data <= 8'h00;
            14'd8323: data <= 8'h00;
            14'd8324: data <= 8'h00;
            14'd8325: data <= 8'h00;
            14'd8326: data <= 8'h0F;
            14'd8327: data <= 8'hFF;
            14'd8328: data <= 8'hFF;
            14'd8329: data <= 8'hFF;
            14'd8330: data <= 8'hFF;
            14'd8331: data <= 8'hFF;
            14'd8332: data <= 8'hFF;
            14'd8333: data <= 8'hFF;
            14'd8334: data <= 8'hFF;
            14'd8335: data <= 8'hFF;
            14'd8336: data <= 8'hFF;
            14'd8337: data <= 8'hC0;
            14'd8338: data <= 8'h1F;
            14'd8339: data <= 8'hFF;
            14'd8340: data <= 8'hFF;
            14'd8341: data <= 8'hFF;
            14'd8342: data <= 8'h8F;
            14'd8343: data <= 8'hFF;
            14'd8344: data <= 8'hFF;
            14'd8345: data <= 8'hFF;
            14'd8346: data <= 8'hFF;
            14'd8347: data <= 8'hFF;
            14'd8348: data <= 8'hFF;
            14'd8349: data <= 8'hFF;
            14'd8350: data <= 8'hFF;
            14'd8351: data <= 8'hFF;
            14'd8352: data <= 8'hFF;
            14'd8353: data <= 8'hF0;
            14'd8354: data <= 8'h00;
            14'd8355: data <= 8'h00;
            14'd8356: data <= 8'h00;
            14'd8357: data <= 8'h00;
            14'd8358: data <= 8'h00;
            14'd8359: data <= 8'h00;
            14'd8360: data <= 8'h00;
            14'd8361: data <= 8'h00;
            14'd8362: data <= 8'h00;
            14'd8363: data <= 8'h00;
            14'd8364: data <= 8'h00;
            14'd8365: data <= 8'h00;
            14'd8366: data <= 8'h0F;
            14'd8367: data <= 8'hFF;
            14'd8368: data <= 8'hFF;
            14'd8369: data <= 8'hFF;
            14'd8370: data <= 8'hFF;
            14'd8371: data <= 8'hFF;
            14'd8372: data <= 8'hFF;
            14'd8373: data <= 8'hFF;
            14'd8374: data <= 8'hFF;
            14'd8375: data <= 8'hFF;
            14'd8376: data <= 8'hFF;
            14'd8377: data <= 8'hF8;
            14'd8378: data <= 8'h3F;
            14'd8379: data <= 8'hFF;
            14'd8380: data <= 8'hFF;
            14'd8381: data <= 8'hFF;
            14'd8382: data <= 8'h87;
            14'd8383: data <= 8'hFF;
            14'd8384: data <= 8'hFF;
            14'd8385: data <= 8'hFF;
            14'd8386: data <= 8'hFF;
            14'd8387: data <= 8'hFF;
            14'd8388: data <= 8'hFF;
            14'd8389: data <= 8'hFF;
            14'd8390: data <= 8'hFF;
            14'd8391: data <= 8'hFF;
            14'd8392: data <= 8'hFF;
            14'd8393: data <= 8'hF0;
            14'd8394: data <= 8'h00;
            14'd8395: data <= 8'h00;
            14'd8396: data <= 8'h00;
            14'd8397: data <= 8'h00;
            14'd8398: data <= 8'h00;
            14'd8399: data <= 8'h00;
            14'd8400: data <= 8'h00;
            14'd8401: data <= 8'h00;
            14'd8402: data <= 8'h00;
            14'd8403: data <= 8'h00;
            14'd8404: data <= 8'h00;
            14'd8405: data <= 8'h00;
            14'd8406: data <= 8'h0F;
            14'd8407: data <= 8'hFF;
            14'd8408: data <= 8'hFF;
            14'd8409: data <= 8'hFF;
            14'd8410: data <= 8'hFF;
            14'd8411: data <= 8'hFF;
            14'd8412: data <= 8'hFF;
            14'd8413: data <= 8'hFF;
            14'd8414: data <= 8'hFF;
            14'd8415: data <= 8'hFF;
            14'd8416: data <= 8'hFF;
            14'd8417: data <= 8'hF8;
            14'd8418: data <= 8'h3F;
            14'd8419: data <= 8'hFF;
            14'd8420: data <= 8'hFF;
            14'd8421: data <= 8'hFF;
            14'd8422: data <= 8'hC7;
            14'd8423: data <= 8'hFF;
            14'd8424: data <= 8'hFF;
            14'd8425: data <= 8'hFF;
            14'd8426: data <= 8'hFF;
            14'd8427: data <= 8'hFF;
            14'd8428: data <= 8'hFF;
            14'd8429: data <= 8'hFF;
            14'd8430: data <= 8'hFF;
            14'd8431: data <= 8'hFF;
            14'd8432: data <= 8'hFF;
            14'd8433: data <= 8'hF0;
            14'd8434: data <= 8'h00;
            14'd8435: data <= 8'h00;
            14'd8436: data <= 8'h00;
            14'd8437: data <= 8'h00;
            14'd8438: data <= 8'h00;
            14'd8439: data <= 8'h00;
            14'd8440: data <= 8'h00;
            14'd8441: data <= 8'h00;
            14'd8442: data <= 8'h00;
            14'd8443: data <= 8'h00;
            14'd8444: data <= 8'h00;
            14'd8445: data <= 8'h00;
            14'd8446: data <= 8'h0F;
            14'd8447: data <= 8'hFF;
            14'd8448: data <= 8'hFF;
            14'd8449: data <= 8'hFF;
            14'd8450: data <= 8'hFF;
            14'd8451: data <= 8'hFF;
            14'd8452: data <= 8'hFF;
            14'd8453: data <= 8'hFF;
            14'd8454: data <= 8'hFF;
            14'd8455: data <= 8'hFF;
            14'd8456: data <= 8'hFF;
            14'd8457: data <= 8'hF8;
            14'd8458: data <= 8'h3F;
            14'd8459: data <= 8'hFF;
            14'd8460: data <= 8'hFF;
            14'd8461: data <= 8'hFF;
            14'd8462: data <= 8'hC4;
            14'd8463: data <= 8'h7F;
            14'd8464: data <= 8'hF1;
            14'd8465: data <= 8'hFF;
            14'd8466: data <= 8'hFF;
            14'd8467: data <= 8'hFF;
            14'd8468: data <= 8'hFF;
            14'd8469: data <= 8'hFF;
            14'd8470: data <= 8'hFF;
            14'd8471: data <= 8'hFF;
            14'd8472: data <= 8'hFF;
            14'd8473: data <= 8'hF0;
            14'd8474: data <= 8'h00;
            14'd8475: data <= 8'h00;
            14'd8476: data <= 8'h00;
            14'd8477: data <= 8'h00;
            14'd8478: data <= 8'h00;
            14'd8479: data <= 8'h00;
            14'd8480: data <= 8'h00;
            14'd8481: data <= 8'h00;
            14'd8482: data <= 8'h00;
            14'd8483: data <= 8'h00;
            14'd8484: data <= 8'h00;
            14'd8485: data <= 8'h00;
            14'd8486: data <= 8'h0F;
            14'd8487: data <= 8'hFF;
            14'd8488: data <= 8'hFF;
            14'd8489: data <= 8'hFF;
            14'd8490: data <= 8'hFF;
            14'd8491: data <= 8'hFF;
            14'd8492: data <= 8'hFF;
            14'd8493: data <= 8'hFF;
            14'd8494: data <= 8'hFF;
            14'd8495: data <= 8'hFF;
            14'd8496: data <= 8'hFF;
            14'd8497: data <= 8'h60;
            14'd8498: data <= 8'h00;
            14'd8499: data <= 8'hFF;
            14'd8500: data <= 8'hFF;
            14'd8501: data <= 8'hFF;
            14'd8502: data <= 8'hC0;
            14'd8503: data <= 8'h7F;
            14'd8504: data <= 8'hF0;
            14'd8505: data <= 8'hFF;
            14'd8506: data <= 8'hFF;
            14'd8507: data <= 8'hFF;
            14'd8508: data <= 8'hFF;
            14'd8509: data <= 8'hFF;
            14'd8510: data <= 8'hFF;
            14'd8511: data <= 8'hFF;
            14'd8512: data <= 8'hFF;
            14'd8513: data <= 8'hF0;
            14'd8514: data <= 8'h00;
            14'd8515: data <= 8'h00;
            14'd8516: data <= 8'h00;
            14'd8517: data <= 8'h00;
            14'd8518: data <= 8'h00;
            14'd8519: data <= 8'h00;
            14'd8520: data <= 8'h00;
            14'd8521: data <= 8'h00;
            14'd8522: data <= 8'h00;
            14'd8523: data <= 8'h00;
            14'd8524: data <= 8'h00;
            14'd8525: data <= 8'h00;
            14'd8526: data <= 8'h0F;
            14'd8527: data <= 8'hFF;
            14'd8528: data <= 8'hFF;
            14'd8529: data <= 8'hFF;
            14'd8530: data <= 8'hFF;
            14'd8531: data <= 8'hFF;
            14'd8532: data <= 8'hFF;
            14'd8533: data <= 8'hFF;
            14'd8534: data <= 8'hFF;
            14'd8535: data <= 8'hFF;
            14'd8536: data <= 8'hF0;
            14'd8537: data <= 8'h00;
            14'd8538: data <= 8'h00;
            14'd8539: data <= 8'h1F;
            14'd8540: data <= 8'hFF;
            14'd8541: data <= 8'hFF;
            14'd8542: data <= 8'hE0;
            14'd8543: data <= 8'h7F;
            14'd8544: data <= 8'hF1;
            14'd8545: data <= 8'hFF;
            14'd8546: data <= 8'hFF;
            14'd8547: data <= 8'hFF;
            14'd8548: data <= 8'hFF;
            14'd8549: data <= 8'hFF;
            14'd8550: data <= 8'hFF;
            14'd8551: data <= 8'hFF;
            14'd8552: data <= 8'hFF;
            14'd8553: data <= 8'hF0;
            14'd8554: data <= 8'h00;
            14'd8555: data <= 8'h00;
            14'd8556: data <= 8'h00;
            14'd8557: data <= 8'h00;
            14'd8558: data <= 8'h00;
            14'd8559: data <= 8'h00;
            14'd8560: data <= 8'h00;
            14'd8561: data <= 8'h00;
            14'd8562: data <= 8'h00;
            14'd8563: data <= 8'h00;
            14'd8564: data <= 8'h00;
            14'd8565: data <= 8'h00;
            14'd8566: data <= 8'h0F;
            14'd8567: data <= 8'hFF;
            14'd8568: data <= 8'hFF;
            14'd8569: data <= 8'hFF;
            14'd8570: data <= 8'hFF;
            14'd8571: data <= 8'hFF;
            14'd8572: data <= 8'hFF;
            14'd8573: data <= 8'hFF;
            14'd8574: data <= 8'hFF;
            14'd8575: data <= 8'hFF;
            14'd8576: data <= 8'hE0;
            14'd8577: data <= 8'h00;
            14'd8578: data <= 8'h00;
            14'd8579: data <= 8'h1F;
            14'd8580: data <= 8'hFF;
            14'd8581: data <= 8'hFF;
            14'd8582: data <= 8'hE0;
            14'd8583: data <= 8'h7F;
            14'd8584: data <= 8'hF9;
            14'd8585: data <= 8'hFF;
            14'd8586: data <= 8'hFF;
            14'd8587: data <= 8'hFF;
            14'd8588: data <= 8'hFF;
            14'd8589: data <= 8'hFF;
            14'd8590: data <= 8'hFF;
            14'd8591: data <= 8'hFF;
            14'd8592: data <= 8'hFF;
            14'd8593: data <= 8'hF0;
            14'd8594: data <= 8'h00;
            14'd8595: data <= 8'h00;
            14'd8596: data <= 8'h00;
            14'd8597: data <= 8'h00;
            14'd8598: data <= 8'h00;
            14'd8599: data <= 8'h00;
            14'd8600: data <= 8'h00;
            14'd8601: data <= 8'h00;
            14'd8602: data <= 8'h00;
            14'd8603: data <= 8'h00;
            14'd8604: data <= 8'h00;
            14'd8605: data <= 8'h00;
            14'd8606: data <= 8'h0F;
            14'd8607: data <= 8'hFF;
            14'd8608: data <= 8'hFF;
            14'd8609: data <= 8'hFF;
            14'd8610: data <= 8'hFF;
            14'd8611: data <= 8'hFF;
            14'd8612: data <= 8'hFF;
            14'd8613: data <= 8'hFF;
            14'd8614: data <= 8'hFF;
            14'd8615: data <= 8'hFF;
            14'd8616: data <= 8'hF0;
            14'd8617: data <= 8'h00;
            14'd8618: data <= 8'h00;
            14'd8619: data <= 8'h1F;
            14'd8620: data <= 8'hFF;
            14'd8621: data <= 8'hFF;
            14'd8622: data <= 8'hF0;
            14'd8623: data <= 8'hFF;
            14'd8624: data <= 8'hFF;
            14'd8625: data <= 8'hFF;
            14'd8626: data <= 8'hFF;
            14'd8627: data <= 8'h7F;
            14'd8628: data <= 8'hFF;
            14'd8629: data <= 8'hFF;
            14'd8630: data <= 8'hFF;
            14'd8631: data <= 8'hFF;
            14'd8632: data <= 8'hFF;
            14'd8633: data <= 8'hF0;
            14'd8634: data <= 8'h00;
            14'd8635: data <= 8'h00;
            14'd8636: data <= 8'h00;
            14'd8637: data <= 8'h00;
            14'd8638: data <= 8'h00;
            14'd8639: data <= 8'h00;
            14'd8640: data <= 8'h00;
            14'd8641: data <= 8'h00;
            14'd8642: data <= 8'h00;
            14'd8643: data <= 8'h00;
            14'd8644: data <= 8'h00;
            14'd8645: data <= 8'h00;
            14'd8646: data <= 8'h0F;
            14'd8647: data <= 8'hFF;
            14'd8648: data <= 8'hFF;
            14'd8649: data <= 8'hFF;
            14'd8650: data <= 8'hFF;
            14'd8651: data <= 8'hFF;
            14'd8652: data <= 8'hFF;
            14'd8653: data <= 8'hFF;
            14'd8654: data <= 8'hFF;
            14'd8655: data <= 8'hFF;
            14'd8656: data <= 8'hF8;
            14'd8657: data <= 8'hFF;
            14'd8658: data <= 8'hFF;
            14'd8659: data <= 8'hFF;
            14'd8660: data <= 8'hFF;
            14'd8661: data <= 8'hFF;
            14'd8662: data <= 8'hDE;
            14'd8663: data <= 8'hFF;
            14'd8664: data <= 8'hFF;
            14'd8665: data <= 8'hFF;
            14'd8666: data <= 8'hFF;
            14'd8667: data <= 8'hFF;
            14'd8668: data <= 8'hFF;
            14'd8669: data <= 8'hFF;
            14'd8670: data <= 8'hFF;
            14'd8671: data <= 8'hFF;
            14'd8672: data <= 8'hFF;
            14'd8673: data <= 8'hF0;
            14'd8674: data <= 8'h00;
            14'd8675: data <= 8'h00;
            14'd8676: data <= 8'h00;
            14'd8677: data <= 8'h00;
            14'd8678: data <= 8'h00;
            14'd8679: data <= 8'h00;
            14'd8680: data <= 8'h00;
            14'd8681: data <= 8'h00;
            14'd8682: data <= 8'h00;
            14'd8683: data <= 8'h00;
            14'd8684: data <= 8'h00;
            14'd8685: data <= 8'h00;
            14'd8686: data <= 8'h0F;
            14'd8687: data <= 8'hFF;
            14'd8688: data <= 8'hFF;
            14'd8689: data <= 8'hFF;
            14'd8690: data <= 8'hFF;
            14'd8691: data <= 8'hFF;
            14'd8692: data <= 8'hFF;
            14'd8693: data <= 8'hFF;
            14'd8694: data <= 8'hF9;
            14'd8695: data <= 8'hFF;
            14'd8696: data <= 8'hFF;
            14'd8697: data <= 8'hFF;
            14'd8698: data <= 8'hFF;
            14'd8699: data <= 8'hFF;
            14'd8700: data <= 8'hFF;
            14'd8701: data <= 8'hFF;
            14'd8702: data <= 8'hEF;
            14'd8703: data <= 8'hFF;
            14'd8704: data <= 8'hFF;
            14'd8705: data <= 8'hFF;
            14'd8706: data <= 8'hFF;
            14'd8707: data <= 8'hFF;
            14'd8708: data <= 8'hFF;
            14'd8709: data <= 8'hFF;
            14'd8710: data <= 8'hFF;
            14'd8711: data <= 8'hFF;
            14'd8712: data <= 8'hFF;
            14'd8713: data <= 8'hF0;
            14'd8714: data <= 8'h00;
            14'd8715: data <= 8'h00;
            14'd8716: data <= 8'h00;
            14'd8717: data <= 8'h00;
            14'd8718: data <= 8'h00;
            14'd8719: data <= 8'h00;
            14'd8720: data <= 8'h00;
            14'd8721: data <= 8'h00;
            14'd8722: data <= 8'h00;
            14'd8723: data <= 8'h00;
            14'd8724: data <= 8'h00;
            14'd8725: data <= 8'h00;
            14'd8726: data <= 8'h0F;
            14'd8727: data <= 8'hFF;
            14'd8728: data <= 8'hFF;
            14'd8729: data <= 8'hFF;
            14'd8730: data <= 8'hFF;
            14'd8731: data <= 8'hFF;
            14'd8732: data <= 8'hFF;
            14'd8733: data <= 8'hFF;
            14'd8734: data <= 8'hFF;
            14'd8735: data <= 8'hFF;
            14'd8736: data <= 8'hFF;
            14'd8737: data <= 8'hFF;
            14'd8738: data <= 8'hFF;
            14'd8739: data <= 8'hFF;
            14'd8740: data <= 8'hFF;
            14'd8741: data <= 8'hFF;
            14'd8742: data <= 8'hFF;
            14'd8743: data <= 8'hFF;
            14'd8744: data <= 8'hFF;
            14'd8745: data <= 8'hFF;
            14'd8746: data <= 8'hFF;
            14'd8747: data <= 8'hFF;
            14'd8748: data <= 8'hFF;
            14'd8749: data <= 8'hFF;
            14'd8750: data <= 8'hFF;
            14'd8751: data <= 8'hFF;
            14'd8752: data <= 8'hFF;
            14'd8753: data <= 8'hF0;
            14'd8754: data <= 8'h00;
            14'd8755: data <= 8'h00;
            14'd8756: data <= 8'h00;
            14'd8757: data <= 8'h00;
            14'd8758: data <= 8'h00;
            14'd8759: data <= 8'h00;
            14'd8760: data <= 8'h00;
            14'd8761: data <= 8'h00;
            14'd8762: data <= 8'h00;
            14'd8763: data <= 8'h00;
            14'd8764: data <= 8'h00;
            14'd8765: data <= 8'h00;
            14'd8766: data <= 8'h0F;
            14'd8767: data <= 8'hFF;
            14'd8768: data <= 8'hFF;
            14'd8769: data <= 8'hFF;
            14'd8770: data <= 8'hFF;
            14'd8771: data <= 8'hFF;
            14'd8772: data <= 8'hFF;
            14'd8773: data <= 8'hFF;
            14'd8774: data <= 8'hFF;
            14'd8775: data <= 8'hFF;
            14'd8776: data <= 8'hFF;
            14'd8777: data <= 8'hFF;
            14'd8778: data <= 8'hFF;
            14'd8779: data <= 8'hFF;
            14'd8780: data <= 8'hFF;
            14'd8781: data <= 8'hFF;
            14'd8782: data <= 8'hFF;
            14'd8783: data <= 8'hFF;
            14'd8784: data <= 8'hFF;
            14'd8785: data <= 8'hFF;
            14'd8786: data <= 8'hFF;
            14'd8787: data <= 8'hFF;
            14'd8788: data <= 8'hFF;
            14'd8789: data <= 8'hFF;
            14'd8790: data <= 8'hFF;
            14'd8791: data <= 8'hFF;
            14'd8792: data <= 8'hFF;
            14'd8793: data <= 8'hF0;
            14'd8794: data <= 8'h00;
            14'd8795: data <= 8'h00;
            14'd8796: data <= 8'h00;
            14'd8797: data <= 8'h00;
            14'd8798: data <= 8'h00;
            14'd8799: data <= 8'h00;
            14'd8800: data <= 8'h00;
            14'd8801: data <= 8'h00;
            14'd8802: data <= 8'h00;
            14'd8803: data <= 8'h00;
            14'd8804: data <= 8'h00;
            14'd8805: data <= 8'h00;
            14'd8806: data <= 8'h0F;
            14'd8807: data <= 8'hFF;
            14'd8808: data <= 8'hFF;
            14'd8809: data <= 8'hFF;
            14'd8810: data <= 8'hFF;
            14'd8811: data <= 8'hFF;
            14'd8812: data <= 8'hFF;
            14'd8813: data <= 8'hFF;
            14'd8814: data <= 8'hFF;
            14'd8815: data <= 8'hFF;
            14'd8816: data <= 8'hFF;
            14'd8817: data <= 8'hFF;
            14'd8818: data <= 8'hFF;
            14'd8819: data <= 8'hFF;
            14'd8820: data <= 8'hFF;
            14'd8821: data <= 8'hFF;
            14'd8822: data <= 8'hFF;
            14'd8823: data <= 8'hFF;
            14'd8824: data <= 8'hFF;
            14'd8825: data <= 8'hFF;
            14'd8826: data <= 8'hFF;
            14'd8827: data <= 8'hFF;
            14'd8828: data <= 8'hFF;
            14'd8829: data <= 8'hFF;
            14'd8830: data <= 8'hFF;
            14'd8831: data <= 8'hFF;
            14'd8832: data <= 8'hFF;
            14'd8833: data <= 8'hF0;
            14'd8834: data <= 8'h00;
            14'd8835: data <= 8'h00;
            14'd8836: data <= 8'h00;
            14'd8837: data <= 8'h00;
            14'd8838: data <= 8'h00;
            14'd8839: data <= 8'h00;
            14'd8840: data <= 8'h00;
            14'd8841: data <= 8'h00;
            14'd8842: data <= 8'h00;
            14'd8843: data <= 8'h00;
            14'd8844: data <= 8'h00;
            14'd8845: data <= 8'h00;
            14'd8846: data <= 8'h0F;
            14'd8847: data <= 8'hFF;
            14'd8848: data <= 8'hFF;
            14'd8849: data <= 8'hFF;
            14'd8850: data <= 8'hFF;
            14'd8851: data <= 8'hFF;
            14'd8852: data <= 8'hFF;
            14'd8853: data <= 8'hFF;
            14'd8854: data <= 8'hFF;
            14'd8855: data <= 8'hFF;
            14'd8856: data <= 8'hFF;
            14'd8857: data <= 8'hFF;
            14'd8858: data <= 8'hFF;
            14'd8859: data <= 8'hFF;
            14'd8860: data <= 8'hFF;
            14'd8861: data <= 8'hFF;
            14'd8862: data <= 8'hFF;
            14'd8863: data <= 8'hFF;
            14'd8864: data <= 8'hFF;
            14'd8865: data <= 8'hFF;
            14'd8866: data <= 8'hFF;
            14'd8867: data <= 8'hFF;
            14'd8868: data <= 8'hFF;
            14'd8869: data <= 8'hFF;
            14'd8870: data <= 8'hFF;
            14'd8871: data <= 8'hFF;
            14'd8872: data <= 8'hFF;
            14'd8873: data <= 8'hF0;
            14'd8874: data <= 8'h00;
            14'd8875: data <= 8'h00;
            14'd8876: data <= 8'h00;
            14'd8877: data <= 8'h00;
            14'd8878: data <= 8'h00;
            14'd8879: data <= 8'h00;
            14'd8880: data <= 8'h00;
            14'd8881: data <= 8'h00;
            14'd8882: data <= 8'h00;
            14'd8883: data <= 8'h00;
            14'd8884: data <= 8'h00;
            14'd8885: data <= 8'h00;
            14'd8886: data <= 8'h0F;
            14'd8887: data <= 8'hFF;
            14'd8888: data <= 8'hFF;
            14'd8889: data <= 8'hFF;
            14'd8890: data <= 8'hFF;
            14'd8891: data <= 8'hFF;
            14'd8892: data <= 8'hFF;
            14'd8893: data <= 8'hFF;
            14'd8894: data <= 8'hFF;
            14'd8895: data <= 8'hFF;
            14'd8896: data <= 8'hFF;
            14'd8897: data <= 8'hFF;
            14'd8898: data <= 8'hFF;
            14'd8899: data <= 8'hFF;
            14'd8900: data <= 8'hFF;
            14'd8901: data <= 8'hFF;
            14'd8902: data <= 8'hFF;
            14'd8903: data <= 8'hFF;
            14'd8904: data <= 8'hFF;
            14'd8905: data <= 8'hFF;
            14'd8906: data <= 8'hFF;
            14'd8907: data <= 8'hFF;
            14'd8908: data <= 8'hFF;
            14'd8909: data <= 8'hFF;
            14'd8910: data <= 8'hFF;
            14'd8911: data <= 8'hFF;
            14'd8912: data <= 8'hFF;
            14'd8913: data <= 8'hF0;
            14'd8914: data <= 8'h00;
            14'd8915: data <= 8'h00;
            14'd8916: data <= 8'h00;
            14'd8917: data <= 8'h00;
            14'd8918: data <= 8'h00;
            14'd8919: data <= 8'h00;
            14'd8920: data <= 8'h00;
            14'd8921: data <= 8'h00;
            14'd8922: data <= 8'h00;
            14'd8923: data <= 8'h00;
            14'd8924: data <= 8'h00;
            14'd8925: data <= 8'h00;
            14'd8926: data <= 8'h0F;
            14'd8927: data <= 8'hFF;
            14'd8928: data <= 8'hFF;
            14'd8929: data <= 8'hFF;
            14'd8930: data <= 8'hFF;
            14'd8931: data <= 8'hFF;
            14'd8932: data <= 8'hFF;
            14'd8933: data <= 8'hFF;
            14'd8934: data <= 8'hFF;
            14'd8935: data <= 8'hFF;
            14'd8936: data <= 8'hFF;
            14'd8937: data <= 8'hFF;
            14'd8938: data <= 8'hFF;
            14'd8939: data <= 8'hFF;
            14'd8940: data <= 8'hFF;
            14'd8941: data <= 8'hFF;
            14'd8942: data <= 8'hFF;
            14'd8943: data <= 8'hFF;
            14'd8944: data <= 8'hFF;
            14'd8945: data <= 8'hFF;
            14'd8946: data <= 8'hFF;
            14'd8947: data <= 8'hFF;
            14'd8948: data <= 8'hFF;
            14'd8949: data <= 8'hFF;
            14'd8950: data <= 8'hFF;
            14'd8951: data <= 8'hFF;
            14'd8952: data <= 8'hFF;
            14'd8953: data <= 8'hF0;
            14'd8954: data <= 8'h00;
            14'd8955: data <= 8'h00;
            14'd8956: data <= 8'h00;
            14'd8957: data <= 8'h00;
            14'd8958: data <= 8'h00;
            14'd8959: data <= 8'h00;
            14'd8960: data <= 8'h00;
            14'd8961: data <= 8'h00;
            14'd8962: data <= 8'h00;
            14'd8963: data <= 8'h00;
            14'd8964: data <= 8'h00;
            14'd8965: data <= 8'h00;
            14'd8966: data <= 8'h0F;
            14'd8967: data <= 8'hFF;
            14'd8968: data <= 8'hFF;
            14'd8969: data <= 8'hFF;
            14'd8970: data <= 8'hFF;
            14'd8971: data <= 8'hFF;
            14'd8972: data <= 8'hFF;
            14'd8973: data <= 8'hFF;
            14'd8974: data <= 8'hFF;
            14'd8975: data <= 8'hFF;
            14'd8976: data <= 8'hFF;
            14'd8977: data <= 8'hFF;
            14'd8978: data <= 8'hFF;
            14'd8979: data <= 8'hFF;
            14'd8980: data <= 8'hFF;
            14'd8981: data <= 8'hFF;
            14'd8982: data <= 8'hFF;
            14'd8983: data <= 8'hFF;
            14'd8984: data <= 8'hFF;
            14'd8985: data <= 8'hFF;
            14'd8986: data <= 8'hFF;
            14'd8987: data <= 8'hFF;
            14'd8988: data <= 8'hFF;
            14'd8989: data <= 8'hFF;
            14'd8990: data <= 8'hFF;
            14'd8991: data <= 8'hFF;
            14'd8992: data <= 8'hFF;
            14'd8993: data <= 8'hF0;
            14'd8994: data <= 8'h00;
            14'd8995: data <= 8'h00;
            14'd8996: data <= 8'h00;
            14'd8997: data <= 8'h00;
            14'd8998: data <= 8'h00;
            14'd8999: data <= 8'h00;
            14'd9000: data <= 8'h00;
            14'd9001: data <= 8'h00;
            14'd9002: data <= 8'h00;
            14'd9003: data <= 8'h00;
            14'd9004: data <= 8'h00;
            14'd9005: data <= 8'h00;
            14'd9006: data <= 8'h0F;
            14'd9007: data <= 8'hFF;
            14'd9008: data <= 8'hFF;
            14'd9009: data <= 8'hFF;
            14'd9010: data <= 8'hFF;
            14'd9011: data <= 8'hFF;
            14'd9012: data <= 8'hFF;
            14'd9013: data <= 8'hFF;
            14'd9014: data <= 8'hFF;
            14'd9015: data <= 8'hFF;
            14'd9016: data <= 8'hFF;
            14'd9017: data <= 8'hFF;
            14'd9018: data <= 8'hFF;
            14'd9019: data <= 8'hFF;
            14'd9020: data <= 8'hFF;
            14'd9021: data <= 8'hFF;
            14'd9022: data <= 8'hFF;
            14'd9023: data <= 8'hFF;
            14'd9024: data <= 8'hFF;
            14'd9025: data <= 8'hFF;
            14'd9026: data <= 8'hFF;
            14'd9027: data <= 8'hFF;
            14'd9028: data <= 8'hFF;
            14'd9029: data <= 8'hFF;
            14'd9030: data <= 8'hFF;
            14'd9031: data <= 8'hFF;
            14'd9032: data <= 8'hFF;
            14'd9033: data <= 8'hF0;
            14'd9034: data <= 8'h00;
            14'd9035: data <= 8'h00;
            14'd9036: data <= 8'h00;
            14'd9037: data <= 8'h00;
            14'd9038: data <= 8'h00;
            14'd9039: data <= 8'h00;
            14'd9040: data <= 8'h00;
            14'd9041: data <= 8'h00;
            14'd9042: data <= 8'h00;
            14'd9043: data <= 8'h00;
            14'd9044: data <= 8'h00;
            14'd9045: data <= 8'h00;
            14'd9046: data <= 8'h0F;
            14'd9047: data <= 8'hFF;
            14'd9048: data <= 8'hFF;
            14'd9049: data <= 8'hFF;
            14'd9050: data <= 8'hFF;
            14'd9051: data <= 8'hFF;
            14'd9052: data <= 8'hFF;
            14'd9053: data <= 8'hFF;
            14'd9054: data <= 8'hFF;
            14'd9055: data <= 8'hFF;
            14'd9056: data <= 8'hFF;
            14'd9057: data <= 8'hFF;
            14'd9058: data <= 8'hFF;
            14'd9059: data <= 8'hFF;
            14'd9060: data <= 8'hFF;
            14'd9061: data <= 8'hFF;
            14'd9062: data <= 8'hFF;
            14'd9063: data <= 8'hFF;
            14'd9064: data <= 8'hFF;
            14'd9065: data <= 8'hFF;
            14'd9066: data <= 8'hFF;
            14'd9067: data <= 8'hFF;
            14'd9068: data <= 8'hFF;
            14'd9069: data <= 8'hFF;
            14'd9070: data <= 8'hFF;
            14'd9071: data <= 8'hFF;
            14'd9072: data <= 8'hFF;
            14'd9073: data <= 8'hF0;
            14'd9074: data <= 8'h00;
            14'd9075: data <= 8'h00;
            14'd9076: data <= 8'h00;
            14'd9077: data <= 8'h00;
            14'd9078: data <= 8'h00;
            14'd9079: data <= 8'h00;
            14'd9080: data <= 8'h00;
            14'd9081: data <= 8'h00;
            14'd9082: data <= 8'h00;
            14'd9083: data <= 8'h00;
            14'd9084: data <= 8'h00;
            14'd9085: data <= 8'h00;
            14'd9086: data <= 8'h0F;
            14'd9087: data <= 8'hFF;
            14'd9088: data <= 8'hFF;
            14'd9089: data <= 8'hFF;
            14'd9090: data <= 8'hFF;
            14'd9091: data <= 8'hFF;
            14'd9092: data <= 8'hFF;
            14'd9093: data <= 8'hFF;
            14'd9094: data <= 8'hFF;
            14'd9095: data <= 8'hFF;
            14'd9096: data <= 8'hFF;
            14'd9097: data <= 8'hFF;
            14'd9098: data <= 8'hFF;
            14'd9099: data <= 8'hFF;
            14'd9100: data <= 8'hFF;
            14'd9101: data <= 8'hF7;
            14'd9102: data <= 8'hFF;
            14'd9103: data <= 8'hFF;
            14'd9104: data <= 8'hFF;
            14'd9105: data <= 8'hFF;
            14'd9106: data <= 8'hFF;
            14'd9107: data <= 8'hFF;
            14'd9108: data <= 8'hFF;
            14'd9109: data <= 8'hFF;
            14'd9110: data <= 8'hFF;
            14'd9111: data <= 8'hFF;
            14'd9112: data <= 8'hFF;
            14'd9113: data <= 8'hF0;
            14'd9114: data <= 8'h00;
            14'd9115: data <= 8'h00;
            14'd9116: data <= 8'h00;
            14'd9117: data <= 8'h00;
            14'd9118: data <= 8'h00;
            14'd9119: data <= 8'h00;
            14'd9120: data <= 8'h00;
            14'd9121: data <= 8'h00;
            14'd9122: data <= 8'h00;
            14'd9123: data <= 8'h00;
            14'd9124: data <= 8'h00;
            14'd9125: data <= 8'h00;
            14'd9126: data <= 8'h0F;
            14'd9127: data <= 8'hFF;
            14'd9128: data <= 8'hFF;
            14'd9129: data <= 8'hFF;
            14'd9130: data <= 8'hFF;
            14'd9131: data <= 8'hFF;
            14'd9132: data <= 8'hFF;
            14'd9133: data <= 8'hFF;
            14'd9134: data <= 8'hFF;
            14'd9135: data <= 8'hFF;
            14'd9136: data <= 8'hFF;
            14'd9137: data <= 8'hFF;
            14'd9138: data <= 8'hFF;
            14'd9139: data <= 8'hFF;
            14'd9140: data <= 8'hFF;
            14'd9141: data <= 8'hFF;
            14'd9142: data <= 8'hFF;
            14'd9143: data <= 8'hFF;
            14'd9144: data <= 8'hFF;
            14'd9145: data <= 8'h7F;
            14'd9146: data <= 8'hFF;
            14'd9147: data <= 8'hFF;
            14'd9148: data <= 8'hFF;
            14'd9149: data <= 8'hFF;
            14'd9150: data <= 8'hFF;
            14'd9151: data <= 8'hFF;
            14'd9152: data <= 8'hFF;
            14'd9153: data <= 8'hF0;
            14'd9154: data <= 8'h00;
            14'd9155: data <= 8'h00;
            14'd9156: data <= 8'h00;
            14'd9157: data <= 8'h00;
            14'd9158: data <= 8'h00;
            14'd9159: data <= 8'h00;
            14'd9160: data <= 8'h00;
            14'd9161: data <= 8'h00;
            14'd9162: data <= 8'h00;
            14'd9163: data <= 8'h00;
            14'd9164: data <= 8'h00;
            14'd9165: data <= 8'h00;
            14'd9166: data <= 8'h0F;
            14'd9167: data <= 8'hFF;
            14'd9168: data <= 8'hFF;
            14'd9169: data <= 8'hFF;
            14'd9170: data <= 8'hFF;
            14'd9171: data <= 8'hFF;
            14'd9172: data <= 8'hFF;
            14'd9173: data <= 8'hFF;
            14'd9174: data <= 8'hFF;
            14'd9175: data <= 8'hFF;
            14'd9176: data <= 8'hFF;
            14'd9177: data <= 8'hFF;
            14'd9178: data <= 8'hFF;
            14'd9179: data <= 8'hFF;
            14'd9180: data <= 8'hFF;
            14'd9181: data <= 8'hFF;
            14'd9182: data <= 8'hFF;
            14'd9183: data <= 8'hFF;
            14'd9184: data <= 8'hFF;
            14'd9185: data <= 8'hFF;
            14'd9186: data <= 8'hFF;
            14'd9187: data <= 8'hFF;
            14'd9188: data <= 8'hFF;
            14'd9189: data <= 8'hFF;
            14'd9190: data <= 8'hFF;
            14'd9191: data <= 8'hFF;
            14'd9192: data <= 8'hFF;
            14'd9193: data <= 8'hF0;
            14'd9194: data <= 8'h00;
            14'd9195: data <= 8'h00;
            14'd9196: data <= 8'h00;
            14'd9197: data <= 8'h00;
            14'd9198: data <= 8'h00;
            14'd9199: data <= 8'h00;
            14'd9200: data <= 8'h00;
            14'd9201: data <= 8'h00;
            14'd9202: data <= 8'h00;
            14'd9203: data <= 8'h00;
            14'd9204: data <= 8'h00;
            14'd9205: data <= 8'h00;
            14'd9206: data <= 8'h0F;
            14'd9207: data <= 8'hFF;
            14'd9208: data <= 8'hFF;
            14'd9209: data <= 8'hFF;
            14'd9210: data <= 8'hFF;
            14'd9211: data <= 8'hFF;
            14'd9212: data <= 8'hFF;
            14'd9213: data <= 8'hFF;
            14'd9214: data <= 8'hFF;
            14'd9215: data <= 8'hFF;
            14'd9216: data <= 8'hFF;
            14'd9217: data <= 8'hFF;
            14'd9218: data <= 8'hFF;
            14'd9219: data <= 8'hFF;
            14'd9220: data <= 8'hFF;
            14'd9221: data <= 8'hFF;
            14'd9222: data <= 8'hFF;
            14'd9223: data <= 8'hFF;
            14'd9224: data <= 8'hFF;
            14'd9225: data <= 8'hFF;
            14'd9226: data <= 8'hFF;
            14'd9227: data <= 8'hFF;
            14'd9228: data <= 8'hFF;
            14'd9229: data <= 8'hFF;
            14'd9230: data <= 8'hFF;
            14'd9231: data <= 8'hFF;
            14'd9232: data <= 8'hFF;
            14'd9233: data <= 8'hF0;
            14'd9234: data <= 8'h00;
            14'd9235: data <= 8'h00;
            14'd9236: data <= 8'h00;
            14'd9237: data <= 8'h00;
            14'd9238: data <= 8'h00;
            14'd9239: data <= 8'h00;
            14'd9240: data <= 8'h00;
            14'd9241: data <= 8'h00;
            14'd9242: data <= 8'h00;
            14'd9243: data <= 8'h00;
            14'd9244: data <= 8'h00;
            14'd9245: data <= 8'h00;
            14'd9246: data <= 8'h0F;
            14'd9247: data <= 8'hFF;
            14'd9248: data <= 8'hFF;
            14'd9249: data <= 8'hFF;
            14'd9250: data <= 8'hFF;
            14'd9251: data <= 8'hFF;
            14'd9252: data <= 8'hFF;
            14'd9253: data <= 8'hFF;
            14'd9254: data <= 8'hFB;
            14'd9255: data <= 8'hFF;
            14'd9256: data <= 8'hFF;
            14'd9257: data <= 8'hFF;
            14'd9258: data <= 8'hFF;
            14'd9259: data <= 8'hFF;
            14'd9260: data <= 8'hFF;
            14'd9261: data <= 8'hFF;
            14'd9262: data <= 8'hFF;
            14'd9263: data <= 8'hFF;
            14'd9264: data <= 8'hFF;
            14'd9265: data <= 8'hFF;
            14'd9266: data <= 8'hFF;
            14'd9267: data <= 8'hFF;
            14'd9268: data <= 8'hFF;
            14'd9269: data <= 8'hFF;
            14'd9270: data <= 8'hFF;
            14'd9271: data <= 8'hFF;
            14'd9272: data <= 8'hFF;
            14'd9273: data <= 8'hF0;
            14'd9274: data <= 8'h00;
            14'd9275: data <= 8'h00;
            14'd9276: data <= 8'h00;
            14'd9277: data <= 8'h00;
            14'd9278: data <= 8'h00;
            14'd9279: data <= 8'h00;
            14'd9280: data <= 8'h00;
            14'd9281: data <= 8'h00;
            14'd9282: data <= 8'h00;
            14'd9283: data <= 8'h00;
            14'd9284: data <= 8'h00;
            14'd9285: data <= 8'h00;
            14'd9286: data <= 8'h0F;
            14'd9287: data <= 8'hFF;
            14'd9288: data <= 8'hFF;
            14'd9289: data <= 8'hFF;
            14'd9290: data <= 8'hFF;
            14'd9291: data <= 8'hFF;
            14'd9292: data <= 8'hFF;
            14'd9293: data <= 8'hFF;
            14'd9294: data <= 8'hFF;
            14'd9295: data <= 8'hFF;
            14'd9296: data <= 8'hFF;
            14'd9297: data <= 8'hFF;
            14'd9298: data <= 8'hFF;
            14'd9299: data <= 8'hFF;
            14'd9300: data <= 8'hFF;
            14'd9301: data <= 8'hFF;
            14'd9302: data <= 8'hFF;
            14'd9303: data <= 8'hFF;
            14'd9304: data <= 8'hFF;
            14'd9305: data <= 8'hFF;
            14'd9306: data <= 8'hFF;
            14'd9307: data <= 8'hFF;
            14'd9308: data <= 8'hFF;
            14'd9309: data <= 8'hFF;
            14'd9310: data <= 8'hFF;
            14'd9311: data <= 8'hFF;
            14'd9312: data <= 8'hFF;
            14'd9313: data <= 8'hF0;
            14'd9314: data <= 8'h00;
            14'd9315: data <= 8'h00;
            14'd9316: data <= 8'h00;
            14'd9317: data <= 8'h00;
            14'd9318: data <= 8'h00;
            14'd9319: data <= 8'h00;
            14'd9320: data <= 8'h00;
            14'd9321: data <= 8'h00;
            14'd9322: data <= 8'h00;
            14'd9323: data <= 8'h00;
            14'd9324: data <= 8'h00;
            14'd9325: data <= 8'h00;
            14'd9326: data <= 8'h0F;
            14'd9327: data <= 8'hFF;
            14'd9328: data <= 8'hFF;
            14'd9329: data <= 8'hFF;
            14'd9330: data <= 8'hFF;
            14'd9331: data <= 8'hFF;
            14'd9332: data <= 8'hFF;
            14'd9333: data <= 8'hFF;
            14'd9334: data <= 8'hFF;
            14'd9335: data <= 8'hFF;
            14'd9336: data <= 8'hFF;
            14'd9337: data <= 8'hFF;
            14'd9338: data <= 8'hFF;
            14'd9339: data <= 8'hFF;
            14'd9340: data <= 8'hFF;
            14'd9341: data <= 8'hFF;
            14'd9342: data <= 8'hFF;
            14'd9343: data <= 8'hFF;
            14'd9344: data <= 8'hFF;
            14'd9345: data <= 8'hFF;
            14'd9346: data <= 8'hFF;
            14'd9347: data <= 8'hFF;
            14'd9348: data <= 8'hFF;
            14'd9349: data <= 8'hFF;
            14'd9350: data <= 8'hFF;
            14'd9351: data <= 8'hFF;
            14'd9352: data <= 8'hFF;
            14'd9353: data <= 8'hF0;
            14'd9354: data <= 8'h00;
            14'd9355: data <= 8'h00;
            14'd9356: data <= 8'h00;
            14'd9357: data <= 8'h00;
            14'd9358: data <= 8'h00;
            14'd9359: data <= 8'h00;
            14'd9360: data <= 8'h00;
            14'd9361: data <= 8'h00;
            14'd9362: data <= 8'h00;
            14'd9363: data <= 8'h00;
            14'd9364: data <= 8'h00;
            14'd9365: data <= 8'h00;
            14'd9366: data <= 8'h0F;
            14'd9367: data <= 8'hFF;
            14'd9368: data <= 8'hFF;
            14'd9369: data <= 8'hFF;
            14'd9370: data <= 8'hFF;
            14'd9371: data <= 8'hFF;
            14'd9372: data <= 8'hFF;
            14'd9373: data <= 8'hFF;
            14'd9374: data <= 8'hFF;
            14'd9375: data <= 8'hFF;
            14'd9376: data <= 8'hFF;
            14'd9377: data <= 8'hFF;
            14'd9378: data <= 8'hFF;
            14'd9379: data <= 8'hFF;
            14'd9380: data <= 8'hFF;
            14'd9381: data <= 8'hFF;
            14'd9382: data <= 8'hFF;
            14'd9383: data <= 8'hFF;
            14'd9384: data <= 8'hFF;
            14'd9385: data <= 8'hFF;
            14'd9386: data <= 8'hFF;
            14'd9387: data <= 8'hFF;
            14'd9388: data <= 8'hFF;
            14'd9389: data <= 8'hFF;
            14'd9390: data <= 8'hFF;
            14'd9391: data <= 8'hFF;
            14'd9392: data <= 8'hFF;
            14'd9393: data <= 8'hF0;
            14'd9394: data <= 8'h00;
            14'd9395: data <= 8'h00;
            14'd9396: data <= 8'h00;
            14'd9397: data <= 8'h00;
            14'd9398: data <= 8'h00;
            14'd9399: data <= 8'h00;
            14'd9400: data <= 8'h00;
            14'd9401: data <= 8'h00;
            14'd9402: data <= 8'h00;
            14'd9403: data <= 8'h00;
            14'd9404: data <= 8'h00;
            14'd9405: data <= 8'h00;
            14'd9406: data <= 8'h0F;
            14'd9407: data <= 8'hFF;
            14'd9408: data <= 8'hFF;
            14'd9409: data <= 8'hFF;
            14'd9410: data <= 8'hFF;
            14'd9411: data <= 8'hFF;
            14'd9412: data <= 8'hFF;
            14'd9413: data <= 8'hFF;
            14'd9414: data <= 8'hFF;
            14'd9415: data <= 8'hFF;
            14'd9416: data <= 8'hFF;
            14'd9417: data <= 8'hFF;
            14'd9418: data <= 8'hFF;
            14'd9419: data <= 8'hFF;
            14'd9420: data <= 8'hFF;
            14'd9421: data <= 8'hFF;
            14'd9422: data <= 8'hFF;
            14'd9423: data <= 8'hFF;
            14'd9424: data <= 8'hFF;
            14'd9425: data <= 8'hFF;
            14'd9426: data <= 8'hFF;
            14'd9427: data <= 8'hFF;
            14'd9428: data <= 8'hFF;
            14'd9429: data <= 8'hFF;
            14'd9430: data <= 8'hFF;
            14'd9431: data <= 8'hFF;
            14'd9432: data <= 8'hFF;
            14'd9433: data <= 8'hF0;
            14'd9434: data <= 8'h00;
            14'd9435: data <= 8'h00;
            14'd9436: data <= 8'h00;
            14'd9437: data <= 8'h00;
            14'd9438: data <= 8'h00;
            14'd9439: data <= 8'h00;
            14'd9440: data <= 8'h00;
            14'd9441: data <= 8'h00;
            14'd9442: data <= 8'h00;
            14'd9443: data <= 8'h00;
            14'd9444: data <= 8'h00;
            14'd9445: data <= 8'h00;
            14'd9446: data <= 8'h0F;
            14'd9447: data <= 8'hFF;
            14'd9448: data <= 8'hFF;
            14'd9449: data <= 8'hFF;
            14'd9450: data <= 8'hFF;
            14'd9451: data <= 8'hFF;
            14'd9452: data <= 8'hFF;
            14'd9453: data <= 8'hFF;
            14'd9454: data <= 8'hFF;
            14'd9455: data <= 8'hFF;
            14'd9456: data <= 8'hFF;
            14'd9457: data <= 8'hFF;
            14'd9458: data <= 8'hFF;
            14'd9459: data <= 8'hFF;
            14'd9460: data <= 8'hFF;
            14'd9461: data <= 8'hFF;
            14'd9462: data <= 8'hFF;
            14'd9463: data <= 8'hFF;
            14'd9464: data <= 8'hFF;
            14'd9465: data <= 8'hFF;
            14'd9466: data <= 8'hFF;
            14'd9467: data <= 8'hFF;
            14'd9468: data <= 8'hFF;
            14'd9469: data <= 8'hFF;
            14'd9470: data <= 8'hFF;
            14'd9471: data <= 8'hFF;
            14'd9472: data <= 8'hFF;
            14'd9473: data <= 8'hF0;
            14'd9474: data <= 8'h00;
            14'd9475: data <= 8'h00;
            14'd9476: data <= 8'h00;
            14'd9477: data <= 8'h00;
            14'd9478: data <= 8'h00;
            14'd9479: data <= 8'h00;
            14'd9480: data <= 8'h00;
            14'd9481: data <= 8'h00;
            14'd9482: data <= 8'h00;
            14'd9483: data <= 8'h00;
            14'd9484: data <= 8'h00;
            14'd9485: data <= 8'h00;
            14'd9486: data <= 8'h0F;
            14'd9487: data <= 8'hFF;
            14'd9488: data <= 8'hFF;
            14'd9489: data <= 8'hFF;
            14'd9490: data <= 8'hFF;
            14'd9491: data <= 8'hFF;
            14'd9492: data <= 8'hFF;
            14'd9493: data <= 8'hFF;
            14'd9494: data <= 8'hFF;
            14'd9495: data <= 8'hFF;
            14'd9496: data <= 8'hFF;
            14'd9497: data <= 8'hFF;
            14'd9498: data <= 8'hFF;
            14'd9499: data <= 8'hFF;
            14'd9500: data <= 8'hFF;
            14'd9501: data <= 8'hFF;
            14'd9502: data <= 8'hFF;
            14'd9503: data <= 8'hFF;
            14'd9504: data <= 8'hFF;
            14'd9505: data <= 8'hFF;
            14'd9506: data <= 8'hFF;
            14'd9507: data <= 8'hFF;
            14'd9508: data <= 8'hFF;
            14'd9509: data <= 8'hFF;
            14'd9510: data <= 8'hFF;
            14'd9511: data <= 8'hFF;
            14'd9512: data <= 8'hFF;
            14'd9513: data <= 8'hF0;
            14'd9514: data <= 8'h00;
            14'd9515: data <= 8'h00;
            14'd9516: data <= 8'h00;
            14'd9517: data <= 8'h00;
            14'd9518: data <= 8'h00;
            14'd9519: data <= 8'h00;
            14'd9520: data <= 8'h00;
            14'd9521: data <= 8'h00;
            14'd9522: data <= 8'h00;
            14'd9523: data <= 8'h00;
            14'd9524: data <= 8'h00;
            14'd9525: data <= 8'h00;
            14'd9526: data <= 8'h0F;
            14'd9527: data <= 8'hFF;
            14'd9528: data <= 8'hFF;
            14'd9529: data <= 8'hFF;
            14'd9530: data <= 8'hFF;
            14'd9531: data <= 8'hFF;
            14'd9532: data <= 8'hFF;
            14'd9533: data <= 8'hFF;
            14'd9534: data <= 8'hFF;
            14'd9535: data <= 8'hFF;
            14'd9536: data <= 8'hFF;
            14'd9537: data <= 8'hFF;
            14'd9538: data <= 8'hFF;
            14'd9539: data <= 8'hFF;
            14'd9540: data <= 8'hFF;
            14'd9541: data <= 8'hFF;
            14'd9542: data <= 8'hFF;
            14'd9543: data <= 8'hFF;
            14'd9544: data <= 8'hFF;
            14'd9545: data <= 8'hFF;
            14'd9546: data <= 8'hFF;
            14'd9547: data <= 8'hFF;
            14'd9548: data <= 8'hFF;
            14'd9549: data <= 8'hFF;
            14'd9550: data <= 8'hFF;
            14'd9551: data <= 8'hFF;
            14'd9552: data <= 8'hFF;
            14'd9553: data <= 8'hF0;
            14'd9554: data <= 8'h00;
            14'd9555: data <= 8'h00;
            14'd9556: data <= 8'h00;
            14'd9557: data <= 8'h00;
            14'd9558: data <= 8'h00;
            14'd9559: data <= 8'h00;
            14'd9560: data <= 8'h00;
            14'd9561: data <= 8'h00;
            14'd9562: data <= 8'h00;
            14'd9563: data <= 8'h00;
            14'd9564: data <= 8'h00;
            14'd9565: data <= 8'h00;
            14'd9566: data <= 8'h0F;
            14'd9567: data <= 8'hFF;
            14'd9568: data <= 8'hFF;
            14'd9569: data <= 8'hFF;
            14'd9570: data <= 8'hFF;
            14'd9571: data <= 8'hFF;
            14'd9572: data <= 8'hFF;
            14'd9573: data <= 8'hFF;
            14'd9574: data <= 8'hFF;
            14'd9575: data <= 8'hFF;
            14'd9576: data <= 8'hFF;
            14'd9577: data <= 8'hFF;
            14'd9578: data <= 8'hFF;
            14'd9579: data <= 8'hFF;
            14'd9580: data <= 8'hFF;
            14'd9581: data <= 8'hFF;
            14'd9582: data <= 8'hFF;
            14'd9583: data <= 8'hFF;
            14'd9584: data <= 8'hFF;
            14'd9585: data <= 8'hFF;
            14'd9586: data <= 8'hFF;
            14'd9587: data <= 8'hFF;
            14'd9588: data <= 8'hFF;
            14'd9589: data <= 8'hFF;
            14'd9590: data <= 8'hFF;
            14'd9591: data <= 8'hFF;
            14'd9592: data <= 8'hFF;
            14'd9593: data <= 8'hF0;
            14'd9594: data <= 8'h00;
            14'd9595: data <= 8'h00;
            14'd9596: data <= 8'h00;
            14'd9597: data <= 8'h00;
            14'd9598: data <= 8'h00;
            14'd9599: data <= 8'h00;
            default: data <= 8'h00;
        endcase
    end

endmodule
